`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
dZwLswzb6oIQsRpZngon6ZH5D4lDooARbLr6wMiSoyNmV5z98++s3WeWw/qB8/QzLZad8bYSfW+B
hyRTZo12YA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aIzvR0PXf1KfOFoAAxi3iy4SUQBu+kkIIVESs7xYjZYa9FMkIi9XvBy3sZ3qYMh26vuV1rRusqK3
kOCxTT/rW4HR/eLa7w8xM4Rp23eDMx0U9TQlkEvboJ3qusYiep+QlJrs6Z87T5Pt5za1/LDZHGNF
nvWAtfW604gJCWi0wjo=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
iHpC6CVvdesjBNk/rV95F+WVZAKIPEDwYCoYioeUYnsnawp09SfvaYAFl5B8M7YmkdzjBfJRumku
Wn8EUsoL1FUV/h3tO3CDWh113sJoeTg0raPjChL5YoHb20nL4ZFp9rpzfwGOdm42mkj5ft/YmvIE
T2S5OxJUqVTznJGk8Iw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
IijTo3b2yr38aI8ErqZlI2TScKXMvmgBX4JZ+BluZRWzUBByNUDHsGxF1Q+5uHzqYKBvOgrIcFK8
Itm8WKbO+oxxkkSK0w7XeoSefxMN3pMQC5hdQdi43Rco78ZkEggSx4KB1tesb9h+rawHDOVlR1Uo
WLKXsfiS49w0NX9PYFCHinwr3VKZ6WxY8tBK/70xTQaBSIGMvp4ygyG5CbXRk1ocOwEgEe/+dOUa
SS+MTyYmju8qAR0ROyf47GWfyMb1yxv5ErgRpwZqwWH5oZxNbURbuczcB5lnav+PJWM+vq9yn4ZK
l8qMjKfSl2zt899b1Ruwa0/u72Kmu+khr1S4dg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
jSf62o5nW+1mSKZKvZ+VxHeCyyNyNCFaVg0MvKdChvOUGyQLgkaqU8dnq9uzDb9brR8MJxZUNnKn
qqXk3k8Gg2r6G0OJNauMh0A7i+x6YPrJYGGII0RyJ0Zmivsri/ZYK5vkZbOjbZkFjHMb9NNXO9f4
LWGE4ln31sDH58U+TOjiqU6Lwa6OxFmMbHmtIjp4iGWwz2263Tfooz7Rf+opvKVu1yfAPtvyXmUo
FAH9P89U292vHW1QA5TtiVTbhdlgOffbyo2/08x0NLH9e0ZM2d96ni669FmeQTYmOutdw/priMj0
7LsOqfvZ/Z0CxT6SMNze9rWCbQ1N3xhUKYptBg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
pL5E0yc+hPF1Lm5RULUIN3nG4cfcDogfXCTgM65aZfAhkqAkt+15bSgVWTqBhUkRKSlsgS5jia/O
WJy2tOudjG34iDoIfeb5XrU7WZ/CFPp8rmT8h6VkrItsDLmXj9RcQeuDAb+k9NPixwcqgdha8Gq0
jv2vezxYZs7uFdqzfhgPugpj08U9mxLLaEfTqi4eFCme6u2jO6HPtupw/IuZVkGuAEXp7Q5OlG2x
Zj8EnNIcofO0En1WPZIBApPLwDsKLhh6I4JgR/BJJiqtPByo4CqvHeEgnwrUCMKhcWZxCrMJxOwN
x1YV0zU3fhscUYzJfyQpDP8AwZE1zN+u9CG6og==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
K/o2RWPX1jSJgtj1GMXJtlz1Q5R6IjkVyc/ACrJ8ybxU4Rw0rglKuz+bTAQYXGsfukgUnh0daHYa
jn0L0grEPW9vqcVv3XT8+Sq7sxNfCCqYGptoswkBRWlUXY0hpO36ePjsY5dhTPIFkAVpLcvcl6pF
A/I1F97b1X73D/K120TMYo7DNfjaOxL2OTT3hoxKevnNo4BkFaEyt7mZX3CQo4pFF4X2YbVEqioX
1M27QB0wQg8Aq0Lrrb3kLGt3pdGI04re3AvrTaXL4fD4kpnrOpQfyC1S2Pd2UykBlap07vaCjFaE
5Dn2ndJTNkeLKnmYP3t4HANuNSOSkeVIK5TinYoAZORhNGUUjaBrRjM32WSJTsEZnqFWE9TV+dau
tnr+eSHtltS2Aw44SnjmvGixH5nU+d5L3IMkY+0LUPnE9tlS3pDxpyno9mlz7txBzXNqLR2I4zKf
nY2XmExKc+VzpLhGSsQcuaZa/3cX9Jxby1ZIiXOdMwhE0MdPwb9nVpFu1D2mMD0OMhIop1YBAUIS
Q2npUbDggw7RI65acJG3gksPJ72rAofDJUtRU/UM3bkmRFzXU8zW50y+rFYkcCu33Nas66qayYbA
8NTdRmSwmGWDcd1QhUUOfrFd6v/1gyNmw3SKneA2kaUwzupd5rywsdGUcxpOIQop5kqlT8wC+gHF
OnAvaElHv4P8QWHZkhtRlpoSJbPogHr9YqFL8NDIfTskrllmH5hyvhWgB5COL4pIZgqv/cvaIkgZ
r6Of8/NV05AKvb9PQAZ1IyS1v/oxM8+rCINfMDKEKWjErwAeopmFo4wUBBLbPhnvVLBAlnOMwwCg
0nA2kJpHhkQHMlZNYgxqaSJmnStZpJbBuisJeA2akqEYx8QfwXP/UmrovK3md1zKnRRVvA1aaiGz
b8hS+t/LuQFHj8JhB407yMJyFwSNhNxTxcWfIxu+xF6rwRamzAPx4nC9q0/HBUl86gL8xQjSI9r6
ksQYD7XpH6MUf56xIw89B+Za9IwINo79WTHUYWYUU8A5d8ukNyPSG3M0IAsbdTgqSC4ydyOHRnmr
ezI/RjKU6+dF4qjAIme/BPn0qc2vOCvDpeaqPBFiZ7Y9OjcfpK+DYG7L8SkTMM+PUc4dDiDCuer4
VsCvgPkrhgMEtBJ8bJGM89hKT03cUQYKdzu2Cczz/SMI6IqGJwoGtIMYzKvI9Hq6nTYFd4nAQkOe
ASN1AYWzfBgHpKR0dUtAs/gikVCYoJvaQGL5KT6ewvcZGbkOCuf0ONd36e1wXeEPmJ6aIcxlFBdW
T4ojsfR/TYZGP4SCA+qBaRuCHFb0zOY8ihNCOCFbhmxtIQQcSnxb3FPWz/orXXXSzuIzd+pHLlTO
XfHCXmbzXVx5JD4mhxzNMe/NTiMifnQRv6213ZICh1v85zUJmisuoSvz4WDs227ufeqxE3GX2SMn
wQFg0JfIZrOjSG0eHku2W8ei/jU/lJpujjk/wWKleoBFcOKwobtz+xWsr/KdKXP3xSuDhEX7i+zQ
wEzWnSjtQiUAZLZbJP3k2+vVYayaY6KzFsxKxwZ11vZHBfSM50eT291VyieVyMu7VZAVmGpoNfdM
dOnuonCFefmO3zdWW8XJgszn+Xa7LsyD9rl/n/Pqe+86ejax25KwXD7LXS5ceU0eW55fwJg52jK6
C1F2Xubfyw0UdJpy32RMVNU47CC9jNVeAVCJAoX/v7tnl2atfy9OfBMS66nfLQfkkx7G9jzca7zm
xny+faHM+Qc2RWQVxIwJBnR/8qvc92vwP+p2h9WiO3IC0UG8bgzGUAtxptiotrmmi9Tf7gCH3no5
5DIOL0xcEqfQMHMC3xrBoW5oIicawMfDRhrTqZ4Cc1C2O4pU9H5ZAowK7BOy6DRf3/DQIcCoM8Ve
hoLNCC5C3stHVOzEVqQIlvIpwXR0GjY4ji08Ie7RraC0s5d6tkMx4ZDiN/gj4MiMCyHaW6Dl5dTu
8HXHMW3wF959EzhzLHWOujbARZBEiRDgNsqzmhPKre+AeDas2IotdX70ddcEllvj2KqcT40trfzB
O19gPBm6NsS4gAikwD59dF5NP55NnXaM7nZddIrOxthGvm8LzKT6dvWIFXIQhkM1NB5+SQ8CO2ZK
AgWyzo3pVxEoorW0R3Covxq2m1ap3x7ipMwAi6qoHKGJgUlgNVgE+unoZbnWue/oQtrIIK6sjwmr
ZhZPac+WV+JzSSeKLJkSwwHbP8WKAtG7py/GTzkpNb5sAEx1LoJa7MQKtp3IwrOrQQDW7nACqoPr
1YmaLxPmMImIYCNl3g2bc+cqGNVz7ZKiCJWRgZrd08Qfdg2VxDgLxp6wMKtDySstJc9Zv5Zgp5TR
Mjec9mz5N1TEgk+/hWzGkSU7+5MIRqPBXRKZTyIvAFiWwnM19HRko7oeCCUsC/4SlMcPRo/Jw4y0
nM0m5hNd/OzVFdz8/3mS3sLzXKAhDpfhCeKHsebyPL6HHXZBB8i/cAXnAyC1Nm6MmSZ/V8GHZcXL
QwiEaLD72As4YWEmTLpfGitxRwOqFrdnM2osRcCAWAai3yT8SDGqfYSR3uj6mmQh9kzX24Z6+FR5
5ugNKBwLhhazyQgiu4VDgEV0E9bwwM2CPeFLrGK4zql0+IXUxWA9XYOGhF9XTKrJrPEhI/EiEwhm
2Niici4HslUSirZ3NNCJ6Fix1qjrno1kSd+gBpekCe2m1tVy+sRBnPcgfp8rl7qAmLRS2TUm4PMu
lS69DqAfz/0tTKiEvdkp6fd8usDYOFFvSUPQtrWDio2nl/guxD+Easq9CrgMJFmgVB8slKCAIgYe
B3+A3Lg1lgRSz0vMnlGl9Sz4xXgL/Kw7LnEIqL79+NIuVMuE3mniIqCzqcCuGcpToRGXeW9cULyz
TS2mz27c5jxYAr6wzTEOWsOIOdRxeX0l0kVGk8JsqjGhWAg/5ar+NmEgYN8+95p1xmqpQnot9wGy
nIQw138KYXFPpNx3jJS13PzqTZyTWseto/7hXUwPwsjKsRlZxJ0XM+ps6XL3pmWBEjKaW4kTZs5j
ZDBRo/twruJ6YuHUbtFE02QyboG6bfvQun1dQ4vJ1CdB8K73+dfLhBhVuzS9yuHGuWM6rn8r+4y2
j/Fj9pWxUf7F69gKjFArFe1HX36WQn2dMJlp9kFMhPmLLcCY4pHG9tnqbDIgX6PkVfRWiHp+dETM
HR2Gh3XaiSenOxGbJXVG+HmFgh+gH2gCuNgUUYyBq1l8KRPfpzGkZpRZ+S2EaHkMgO84rq4rFwtO
YN/H54iE966dp09gXKSCWDt34PRPtN3tBUt4+aZmG15QCz7FMVsgsNcPnl9zA2WceyaUaDURNwfY
TZ9/WTzRUgsyMM4M0JSGnw12riQ7BdkiSVl/eCb6NppDTbsCN0pDq0hoKTlH1RD86ji3xm85YpxP
glyzFiJhh7cmGobpHVOaI9dBhkL9lGzmDH9xMwDdpjbLA1H9IF3WIFk67Khy22I38/TVWlplZJ4H
SrqgmIMXsNh7a4DN1EDLEavYOGNFjfriZ85Nq3R+drRQhNjyNnPklxDIC9VhgtWWsi5pQ2Lkw7NW
SJNrmBzipkt8ndmMdEJio5Asi4PiDjc/PfRyeH8akj5ByChpirSTYVDTqmYTpry+CwNQStc8x606
vvPeKqzn0c/GVL/dhNycKek6Ga2Sp/urCavE9kLx3NL6QQswccrgGO0rNoAOslyv3l1PwyiHl/og
s2MPZHpoStIytq2uuVatCcVn5Mb3eqa5XVl5IPlF3GzvcTT5Aka92pDaKkcHSVALFAL05SAKRwTh
A6Pfc9lW104EID7RJffKV8Gq9ccVgdamrvDb/YrMuR4rt9OfdYYxKPtH/D61VhcGsqQ66cxhhFqs
uL6/ELBytdBQVjgmwPYnRT4z3PpcdZFq0SfxV/k5BU7uzIt25Hw2oi7sMjqF8zx8xv2OZ8T4/FSG
fE8+KYFvfRwY63tZijXS92VkWfXlwZTPuUJLe8JZHkUYdiL4/Ijv6DOuSsEgOzSApFA17GCNuWtw
qki3Ogr3x15SOmHfj1hewvWRfmCKZ/B9c4Ish8GmLT2K7W/uzaq+61YvQam8jI0DKe1ztroL/va3
4OoalMSwZz78bEXYdqa7PRaUySm6vVuPnYwuJvikwk784qaeze96q3PHoNaibdhHVrY+2ndraDlT
lw==
`pragma protect end_protected
