module And(input wire A, B,
	   output wire Y);
   assign Y = A & B;   
endmodule
