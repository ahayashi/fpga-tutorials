`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
OCP9udf96pdCNm0dYKrx/XohP8vvJ9tQpvcqLHaq12Om0pnW2Ig+Ht/7gW3OiDnWmmoL1ulC6OiO
egH12+UhSw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XIsAP0w5qKaJeaO9EKCAPRuIg5cejqDyfMeLt14hWU0ow61kmButV7Y6uA6dKrDKFGRMzdCmxgac
wj+4biaA3FS6oU6asBLMDNSIZtjKYZYKb+0nuqOvwlOw4Yz1k3xbyQvUQHpnev243zk8/c8Sel2t
i+M5WZT8R48xVsyKp0I=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
RYo7a+3IoKwiNqFFQu6DsDjbJFLhzrAor/+tIsyVrG/vDBQk/EpEBgcr+ZXtlylhhMqMy7ZgaeIt
D/CE2lZ4hdz59TvrGLmCEda6MYU8F7gAM0kyqmDVEohG9gSmtbvsmJXjVnrIB3t3F2a8yZEzdRVa
kZgdNrc6UZAbdpuWtzw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
07jSbg76uq/Ky4pZdaGRlh+fUYdpWNseYjApMqn00/wWmtPu0arGAGRFzqyKsUsFpb/4c4Mt/zm8
j2cWn/AuxjGezOa3ceOv2MAn815JriFdHtW7afTxN7LDZVE7QyRrII30l0o+bifm+0cLrLNlVu2p
9FMjejWwZGr0gVCrqn60ytxf56AYDGhZ7M6HNMEN6nUi+BCNI3cgVnZm40LyPfIuhSnl4KTgJDK+
5r07yl9o7TLlcc8MHDhfAD/qHtTRc/zCXt15j2Y7LjAmRnRQWqUSp1mZ60SmL3kWqDMBY6FXWWXE
dRWvxmaggOE1Z5miJ4KlJNG9CqogB+m8qLaE9A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MdKe9TRNjCv96Rt7LRh09EkdSx1oNzcND/XlCb5pt3qBiMqbNa6OvpmmKHmM9fJVoqdVARWcHvP2
GidcffzRrrdeissQybLbWQ65wo365Bg+2OKhFEz3LfqODMjGmU4937VIm/V5UBUkdijehxWLVzoi
lWRPh4T3/9f78eZCk0stCbvKdrhb7T+JI0IY3ZT9Wzep2JFsL4LYk3D1mp/rlkwpd2uADd8fSjtB
ukvE8KwvVketjPpYirRfsSQeKTVLYGq/BsBX9vHRsM9dDu01uJoxp0uzLOsn7xDvDon99E1eRifT
NFiYVhdutShoZrV+6LvP1ycpOcLFZPGk+aba4Q==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
m8R66eZJL4RnmoF4fD6R7KoWYg/o7eOca/Fp8eAXAXxK9eqluz/B8Yrrb8W4N+xUghfWV08NaHdH
TMHBxOUrTk7aFAIrOZ/ytiKL30DCZOuOrMUz8SdprG/pqM2BIvLjLpXgWr8xCWGNNqh+InQS9RjG
DZGkdH2BMSb2AYxFst7Hjp+XeI4mTRHcBR/OVyA/P6o8E/yVgh9CHgVFF9G8DgRl57jL+uq+1ouT
M8IXNEXQx7/sVKAPjL2UYdVsFbPM0TLzutHbvIOKimapE7DMgeFCaQrvyjNCaRAwoKQoVlckCMZF
Mihilj82Aa2Jjecpzl8S2CMUOuwlu2D7U0euCA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15104)
`pragma protect data_block
JqPgEjqUAUNBc9n5AZKVoqZAmBDhN2/RTjCt7kT1uRV1kYCbEVOuh1teIsrrvOCXHfeike3WBSM9
jCGCpG47N4q8sCMLmpNgv0YeXJ3kYWwDIh9GhhTh11+2FFcjz8QsVmBcLZeVoKIHtCGj74acu8MP
r5vWmMdZ5LkZ44Nms+8EChTZ0ShW4oGpm+3Mi7uLPj18uOq8Kg9X47wY5qmSyrg11ZoRdGOHB4v+
XPbW9vd7ksMwOkh3DONgzWGr86EYFM0oBTEAL6jsztvx21YUtRUPshtemV8tYYHSg8IGZbEOGblM
N4rKAnAtGEiBUvwAAxvrw5q9BRX2X2q8mFLL6O5+00+slz/TspeadNir/u6/WX+4ylwEoGOIjfgh
mHRhngaCWPoYYvpY1I4YT3AOf7ZkgOLakFOwQPyGLhEOGggDqyBmsT7Fo/WylXuwVr5lYo8UErIS
FhfSEPT4GL717jOxLrLTAVQNuWTNKfQik6ay4LFBjhviItK3R0vxkbQrNXI33L8RzOpMY+ZUwB7p
Ejdz8v5WoaNUUCc0mwpfqxKIJRH1JAkQb3XJtXrqSwSM6SGTZWxhHtfl4Wdethi7f3xkcq8pZ2GL
1GIC+x7QK1ZoLbgjxTc/7kiWTpEdLfQtMKaGNgjS9uM68ceUoXYBL4D/twDH0I+N4TYfh/sg7y6P
CGz8p+Rgx3PwHKiybP5vCZ5otXdgwsisRwKt1G6HeDlM5iXe06/IqFrPKTj8ht0OYx1mzuW4DiwX
jjY9M7ePoIC7X5OFcmInlI2dSs7y2wkwmgAGPlVNUWJ5I04XDeGAAV8E29RTB/9aCllJRUmDvwxS
3PdelCuOB6tYzEsQv9axFNcEekLoK6OiGJbjG6LSYfmbILi7TMG0AbY4QV66v1iHlaSvq3S3QEpn
J8wPQ2+r6KSUj572VuTH0JpKWgHLFeGfK9Sf1UmG5uv77jAnzzhLGDXf/8A43dGnRtNSEmV+0ow6
V1W3tE/5AHtb9S6yj9FyYtvFecIJt6EBa1b49b7oBQqerGVvxI0ABLeIePDepb8ns2S1iPkDoNXH
n3qXMqiFe5uH8tfyjmkkpdKMPNFEAMdDpbthRTqns7Ejh+lGL1EgQQAsGKHD7PdyUB1y/opB9ODe
IvXC+4hds2TbS8FpNFXT+9iR7EBr58rwP4KHC5HfNODibWAx8WriYQWx22elScT5JkVicrjajvJo
gxL7NSG3hnD/6Y3n8UUEaKwdmRLqHTelZBCY47I+phx0x64jV+slRNxa9gsZPBKNWGIItYYFqlCG
k7YfBXSm/AzcfDnQn+1NStp55HMWIMzEp3ShNTd5QIIKEQP3fMQtx+Zique1jvcp5qxYRGU+BCYb
/FIfKWdeUN35A8tWXDh59BnUsLA6JpTu8y9BP9dYCgmu0Ho39yDkIwBx3hqqY39s0EBgZgyXKCDo
wHYm+ysPaQv7TQUfwR/pbLH/4tg2fk+uov3RHOvzYnKjegqGOewDcU2lLnDSXwXLn4YoEPUC42Ml
tFdREPAvpyB1+K90aSV7ctDyF72mxRemE9eKh1fuEvw++sDKVqXkTJwXiaxNOKPIMwT1tdj9qSeO
bnCy4qSK8g1tAswVAlQegFp1MujyKd5Sb39LfKzo7JNFz8FGUlWyHFADhL64xgeH6nKV1cXFBCZc
qWN08N1DDVDiJlZsHFy8Nal4ZrK4swnOwq6NzmAzwpeYeCwe3iAyh/tYoWdibNig2rALVYGmx1Cy
+4HBCUEf7mXwdDREFVBg8QJ7O4/n3XiaZdrK9ctMg6oBouEUU8kmC0k5GUTVVJAMZma9E7Rs/9tO
CjA+KCHAAYxVFtkz/xAfZVo5pWeoCqzB21odtdmudysukpd3Fue1W3rXc2d0R46blo0gLQNWE+O1
rO39BMKH0ge//DYA1vqLIFhAs0lUDs4Hca31meVGEhAvUBsC0UW+Zrob48VmAm+MyL21GgTRv+0R
xfNLz8uNCT5YFflQN8AXURI/MdIlSY15zLTf+5TZCeIjll35V4VXAcQnQGhAmOFaMNxOW0w+vCBT
4bTu5RIwfovHkh8ffaNSZO5PaSt3ES2wkdGN7R/hKuXg+YARah0/4JNmHuL6F+sKx3F/8d9z04N4
iuEr2LoAbZg0+Y7sXJZQpLlj4ER3lg4VgKINJjug6HiEPoMGyWZjNorlmzhuJo/q+mZ96vs7bmLY
CecCXlz6SsRy4GLsgm1PNyalIwXNs+a4sDh1sl6bZxHhDymXW5OpBiab+NrXtSmE4aPfgcHpPbFL
hb8dVkKmUypHg2ReB4z8/Vz8HXPGl2W72h4s2MRk1ZpHHIVWICO0AOryZ9040dXE3y25w3azwYgH
BgraMV6y5/OBrZ7EDLLDTdKlnurAleik1QURgtGn19tNcqDrwnx6X4J0lpUxrBORKUtDy+DFQstd
ImFhNqBcn/zI3siA2nK3MAcCSznUMeosLRTnu7do2arn5/uS6H+lmJUo1MORCgwam0rNpUoDePnY
6bD3I+vVrkm9AbmBGzcLYSNNnsoxAvDCIaQEOv4lZ1u83+c0TF74bCsGoxsonGYoQQNJ5HFFBD9b
CswYXsvPQrVSvoW8wxa7ikMtISA5MY0rqh6rpMKvr6qHnAER3Ig8vMdBld29GKQyc+6V29DNw+vj
5XOyu25s0lo59yo54bx7A1x5FG7+qYFZu23ynNvInQEQCTIZoqU7sWN1cGICQCfoAB5VYfxwpPiE
jkS5fi7G9q9jsT6mLCSnqcguEgrkvNXghqPFmXVOPFlhkExSkjd3GIIpaCLjuQtp46c8uX4LH8GV
JP/wQ1sCCe2JVNNNAdX/r2k+t8IHLdFcs0yxzHE5LzWq5oFomYWjY2cFbp70YhkUbrfoWn9hC9we
yrFwTlXZxkbY+cumpdBMCsYn3m6ZP0FpA4h7SwaHRG4LC73rc0yioQWyhQf/F1WvIxMwbrLw62Bz
da1jWQAtHSkD8lxaQ//+kfGwCOepoXaaZIhsp6HhdR28o4dBGUpo/+6Y/OSWED3LqZqKHWSk0s5M
kiWs7G0JG1BwbWlfZAeZyjff5Mh+wCFO08nKISWU0ifuTIakqEhTzXIm9Y2ZsJbd4iOrLoyOMNpe
DIvIdxzaijt71TeImX9hqjPW9tl/o2TnVE2ZdRAZljyS/rd82k0BZGylpxtJyJKVNJweFJiXbWrs
YKdk2/AKwGQJLofkdJzaj2VUv7OrLafwPpsgEnKSfrr079/2uYs8jZr15yPo8sYWpHkhBJYMlOTf
z7qGUfUa88I16nXeeuKTlCyWeioqOyCKvXeXGJ2wWrP8JSeEHmy/meXBWUsXVhV3hYpLp4rCQJeQ
svDET1l7QWSUooPGYvJ29cG2FwhEOFxzyMo1ncndv1iM63UtABf9wLXwxdpAkIt0UP9qXQvsDeif
8BlZEqmpvNjvOUrYB/kLFg0R16bYnOeq8kHqAWtkbRm3egWUiKlUOjoqf44/sBJVxGvFS3OlgFl5
heQve9jYc6X+NUAni1/fObiY1SkE9w3Z2hU7bV35ktmCwJ7Jz3M5x8lYk3E61OP3L6vU/NAq4YNj
elkObjp9QInbtCqit/zIX3Oyw4WFzIYgaSE4NkddHruN7JWGBTT89xf4TumN0nXkZXoZHJGpj5Yc
/VjwoxQmzLsivXAnkXt6bUSYxKJdhfGXgRIEw16LvrQMsfePkP06BQjtknaBvXQR6i+ONKtjybT8
gsaUPqPx1RrEp94dbwLBeS0sGUYT9Kk1G/S72GssBcXrS5DzvFqbwEECJD0vli1OpKd8ll1BWWra
uNWFWY4D5Wi4x47FQU8cZJM+EsOhYQYNYSA0ejb+fQQs/M5T6AnwVTRgZbqsPJ7RdkeqnfMzogir
jKPyxS9+l9rKhFLVcR23IQYAS6OO9MiOt2BDt56rGEveYVVhr0svdzq2F003xwtuCW1gRAYcO2I1
OTpAXh5esE95Z0Y18PToCAgkupUXwzS6dkJX1afyLPxauxk2TmkZ0/0j/4M3xkKF0KoCdW/Bot0x
58JMEys7xzzqsApSZTOJNqsUvIu3iT/CYU/TBWHt0JP6f/gGCVSvYY+JuLVOkM3JZXcspzRUlLXy
6RlM2mjWBjS33ozSfnRVhcLRZQbcfxk207Qj563q07BR618z1Kaya+0eKcXbNNSltMoyVJQkYa+9
w347Ni/EBvWamDpbBMp6FH5NKOM7RvaxWlBHrdSKhDtJscQM00kDoF0qO4M5HqMDy/euzpxQh6ux
+s378gapzmSkR9uCdvfUd+a/ZmR6qADPclRi4GvvEVkSDvXAp55iOM4oOksXNyBH4Xh3xXwrST1F
hJWeXNn7kSBhMjlfOpTrKfArPHp6XOdXuazXPHJEl4mrj+xvNuGHMbtmYLM48UuBfuwxRLl8bVBn
qJVPz4ZAIoqY/ZIEqbkALIz/Qf+cLG2QR9DeatlswWGzeaWJcwPrvrrYbEVHUeeId/Qsk/y8n8V7
UDc+leVrJUdl/7NGNtA0VfdyGHUELEugrCnAePBrZy5w7NCGTRjz2DemziINeGL12OfCAcEyoM6J
lfM9EsIAqN50cLTC8M5bh5bElmV4b6OtWSeMh8BCEL93HgtgRP9zt2uS2RO3oiv2glfIZgtqb6iJ
Gg9bRCDd6D+EvYWmCsopn/jWu3llQjBb+oAC73lV0Qe1/gyc+WIEyLPCH4Icv6+IONhOFMT6lmpj
J81fa1eQaDIN8RF0m9elFF4nXD9VAbUfdg0/HkiOFsx7IUEecF9UyRtxq7sq2ap6FWRQcXBu6elg
P7B3+zAjKBklpPDmhpHuXfjjr50ZMX5lCDVcwxgF/9oaOCYSaSyrnfHIXWpv27z7RlJDPY67Twmv
LRQ6k4V5k1PkyaFrE6xa6nCoVhQihQwXWwQT5B7zojPl1OeAvrUYJEPLooiYZv104oUnQ+RVFyOM
W4WfYXBFWruCvt7WtE085S0JRMmMafW9Ui5uUeE+nhZxPXtkoUlZ+P4QTCuzPqsw/vyLY92sJWRF
45p8YPGiA9ruSKumxY80x8os/vMtymLFjIZK2Gc3dXlANDZ+BwPLqw0Up1mfLLKkAPRSYj0Fl7WX
ae7PpRshzWjHbdUJCkxjSX9dtMLG27hdsYapm3wRaCYXFBjXxQAGrFdxmEM9niaRmpPRsiYteMLk
xwn4pFMK1Nwae67fVFFCUQG+hkX0OBk5gj5oIYVRerSTtguJRb4mmNSSE3Mq2IZb2vahh1BoU4z9
OS5F8BlHRcQbvZkglybkT9G59nWfI6GUr6k747R8xEeu5bZNq89PnTTOlgy3KfGI+uitx0ga0RKZ
lndjpJArR9xyGlb3ZZnIMMyd2EFj2llQpxjCoy/3UHtvNBUiBGlifLzGKrhVVHIpW7luTn/GsyOC
8iHwisWzE0fqS2VY56AOs4eL0v8WFmbrnt6a0zHRxyQNf9XW12TaFOjlBYO++hX0NHZXTuyX4j3q
j3rAqfhN3WKg65bStvjcnb3i9HNhe09jiFa4aTLAkee3rrEqks4Ks09sQAlBiBHB7tzebhS4Eblo
f3OQtmJevYHaN3y2Zg69NpOBQUmCCYTUFSH2v6nJxH4dG1zucIIme/FO+TOGWiYwQNu00Oof0HBE
TjmFwZXx/nu6B5RT7Gpmu9oc5Ha7r4KsU12IsW3EiG6ougphS3Ov5qJknccJkHr0oGA2w9zoArys
XhZoSKJ/wX31tEraxWth3eTfm6GffK8x4YMgIQ/48rDsCx6LDeyLejoj/+G3TspgVnDloErJHLI/
czUqVJ70TzjpWRc+ASNuGY/2/QV7R/2ApmI3WcJD2gAnl24mq51RYemNxXHf30+rPZ7pcRu/pTZ+
41OFY+vCfXqEEZxCpl6JSgI8K8VYX965+Xig2gc2jpwlyYcdqB0kKLRDdRwD4gNJnnmprgD+8D13
cAa501PeKMK9iP7+McjHVZu1v8BjiRn+zD76l1X566Za5QxsUCNALG3vOs+g13PsSxU8LErCkYTq
T1Tj2txXTme/Bf9hbintsOlLv7VZUMZTwl4t23x/llYywSoZLe0NNZ+CmbpqgzkX0ASAOiCHmq+D
GCkTW364btyGjZSWXHlVUcFFI1vf3lK2kxVdWE3PvWg1xMFdvkeb9nLnAmtDFbF21XtEaw6d9+UC
sPyUExzSDp+t2gr01L4KPxoXdbWF8vUXQ4NvvrVwmN7EyTAFkMWwS65hU6arjFUxlXbf2UAPBBIf
DbQPdyj7QfR2p1aVi8vHMYrGVvVBkwmHykBiP48AULtUoq2tmAisnu/ik+JnQO6q2c7gt9DcSfId
o/FpHWzSxjltcUPCEIU+IA80gvp7HWMTiO+kfUmvkrid9iwSdiYRlRpWzcFh1B0+W0OzNwNuGzfN
s98WCJq9X8CZuVGKIeTGYv5xQch9DLoLE4+0b2a1L/+jliCdd8PRLRtsyeX6k6WoCCFe2W4SJ48I
EZtyEYxsWiVDX596oY5PBA8BgrpdIq2RVWHCgnZKylOEbezixxbpHzF17WIdK8HGzh5C1qhIHj0Y
I1b5HOKFmoK07Fp+ieU4SIUuSxbDRvV/p8EMI8F7nm+4CfFAShXHSm/zwcixzfKm6bqb1dLRJEX3
xeX0jYw1Cz/yCe1BR31Y0YgEMG92pK7VOeyRV8udzAfLOsZdRg6LMkvfZU5Q6Y6br767v2MZDqjd
xERC5aPgx7jyZ2NsvWj3OACI8Dnqx6sq54gMXKb0F7POGtckPrm111YRbnAESRRkMTKvVw1PwbNq
T0VLKekBgDn9DxJPrlaft5UYWzGvkkA6Cn82i9u+yCmllVUMc15WMETTtDLfqMcKTuKrHBu29ziM
7YtgKBd9Hy1MSiahTe4EBOePL5NbYnpGZ+9MJNBo1jvaUQGQ0PSC6Fk8g7zihkYzUpkMTHwuAAy0
zwpr1Xi2l125kM9sczG8uNOCGRnQaLZtQSIWinA5ftI6zJuoxTWFOawCvJFQVTupnARo+y4T3jYb
9wjoUcEh0TWuabH0uQ5Oe0yHRCyDYtW+TIPLtbHmk+XG+OhW6993NwwE1Dwp+Q/zuGpHM1yBcgsO
/ky2V0UXf1yJCdPrTQgiKqb8WVKRa/u/+JCwFoSCPhfETDA1NdnUpuv93svwSXksB97Fq0VgE2JR
rG0VKTyRk1P40P1lDsOYC9otBBmORB1vnv3tqCNqsvM3Z2DzqIMHFJ6oWgH0s34cQCxjijGgFJvi
3ACEov+ByiUoZjDKk/h6GsmzG7QivGL04JQJhIybEMFUdQe6Eq9567arbmRI9qlNdioo+7nijg9u
+GWkbRsti06bzZPK8hYmgpczoQ+JCGlUKY7/tIe9EJsc6+tQkqFrIdlWYSnynDKrSReIjlVhSgza
LUnQxJxv3kGpzW8QanOnAF/Sh+k/Ky0z3kym+PplAemO99hNIxcVWb4JUIxQY362cWEO532T45lL
markokM/pOuSbeFjIbtpJW5nAbvZrR2/01QkW5t9pIpWoho467CjgwEQIeT9rvMxG6Wyqxh89UO9
ULvgicrJXMAgzFxdNQTxDtZITzAjCQpCMsVeKjrwGMLclOvuyU8cLw4x+oT3NTweOt2yuhKY2lzw
5IL/P0EGI0bHZu2hJMnzO+cfN/hZm88HWJDntkp2QoUfo6E5IWAymEwWEfb4hUjxZXBLOqR789mG
zShFSYwQHpWmpF1uSWm1kuSqcPYtassUkM4GV8opdiV6MM0j163IFNIETR07raYDfCMWXeuu0YSo
fUDJAu8QC2H/L9KDZzOZ1c18nh5+w5Vqxe6ZyZFZzuVbxFgXU5+1afO1GicbQg6Qw8/JO49BzaE0
Qmgd0rRivV4ETlyRZgjIGSZsgWJJuaKh7DRrEO8tGac+6amOjsUf5Ex7dkyDZiZ7ricOkukD9iD8
YYIVyp7nt9ktVkPQJXIVXHQfxy1iIl4HOOrUE9+L0VfkO9L/G5k6lXUtwl1L/X48UjYVH7lZSz35
2q/yFwZETeXoorZ57L4QZ117eGvRFhFWaKcGLYQnVQYzOgJbYsh/E2Q/lrjQ7A57caUhQSDTsOtQ
EolsqV4cCRIqIYPRxb+ealoRk1bcoH1quJYJ64qXa+h0SWZcLtLPWY8lkzNfPrmi4PgraLgPv24H
J26ZM7UgIDOdPCHCdkPnGWVAEQOEuHH9rase1w0K3L6gZNV9V8t5EsCUsnl9JE4kr0Ek429PXPd+
lMXXXMmkqc1NBsGBXXB4GfxIVUZc5smQ+Pifb8cBtgL8alZm9o5s60pFtQg8KIBQhldHb1nkMNPf
2NmGbyEbsj0gYxclrXg3GnRYPr6zI5CEK1bEUQLy3GJSQT3NZ4dbI/AaQcOwWXNxGy/yX2e8mPNl
OdDQC5XaHrzSXQqV/AUkTrQGuPZofAHuWpNV5VVsyTdwnCb6qWG5OnEZovVyRxx7dq5cgWZ4fQqR
9/VEj/cB58NIjxlCRKSFkpVo13yPn0odLU77SipVyLobiKT8hx9l6/MD2RVUbydbVTfOygjlgyc7
YG1RGulZtAMytaXKoYZC1uHpQlj/EiFQCcS+iXi2De0xhC2N9wfl4iVCwuRV3srrbJTuHlr2UPGl
trsYZSFV+WnR9Z8jtU37RsbjPs19KCZ/hr4zp0RthzjbIqPnyrpr6hagbS0HSCmvGKsA3PNHHRWo
ePyFsVtyZY52JntAQQgT/7aXfPD98ePnkU6Eb+snWeihWCOn/Q3g1g7JzyG3NpZkpbhKXEq3hV20
ATSL9cxOzCDkqU2qWHe/DzypfOPOPIjiO7SGSykfXdG8WJbKMYqnhMGs9YmFKQq1Eh3UgSJoHmE5
ee4T2bqIOf2WgdwVbMrWilb0qdnBMlBky5gU2gG01pGr7seiGoUXmeWLNnUp59qTk6NpLHLAYnAH
XncL/n+EewzcROng3EIXwCDHi+yOXxZKYxperFeM8UhCQHD94xRg4WkfO3kNnYLCDarrrfhqi/Ba
DwWspNTw6Suruyx9Nhdt5kVhf2+Nfidd/+alwmZglIouF/r17VJMPAN5PkaWhYptlOH64lw9SlcY
fZFylCfKe3nKn/aohsSwzuDIdiGZhOfDN45CBjNdBhUcG3OlWx9PSqbYUQ/S/ufl9tlj5eMyaNVf
LU4We/n8zZsOiuYInf8pEnoXZJs//GMmW2J1W5SoOCu9Ss0cqRUwKMib819EWbsN4PbPF9eEQz/Y
FNh8o/XXzMQN3yVEfFsNMcghhqqmMnHPTefBS+a9zhS3gzuHvVpx0+BoDASUzGgEGfQNSbJfXAOV
QGSl+GfMMkwQxem2aViY2R7Nj+loj6joDXgED3ERVxuTrsJuvqTkgTiax3qAQgOIsalKwDNahrfr
P6GAAQd0yH/MTVdvRwdaezvBXgQy9I+AC+6XPi1bakRpfn3JBvpQkvjs6mayX9G6vp+z7f1TYTw4
KOrAFPjG28SJR09fI874eHX5wywu3T2+MIzk91Qcp2tc36vhVxqpnV9ou4wbla2oPXqzay3zsiPQ
Swr74Njzn/KMSKMrj3rUVTHkoj9D5+LBupMGiR0wbZJt+JALwbfWJ+wgWeRTavRh1ia60m8CDI1v
TlpOTgFzbRX4bersG2yIH2ILtgvSdgjlvmAB0hT63NsvgxBBjmgaYHj4iCn0UaVchPGoBl30OxxM
BSTMBx+P6XMkCil3S9mDz1BiuNDZJPuYPBPwMnyZ0Yhvj/epWcItw01BcIepjKKY42PRCTxgV/9s
SqLIrrH/E/Y3VHblQJ3RE0GNWogFtBKrj0pODW2JlLRZzt+iFkndQO7VYu9CEBZhuvsiy09DNgmm
6AmuAktcLgd5yxpiv+tR+K7utJB/68ruSeEili/U3JT1PT9o33i1dMkLnR87VtI6MFZd1Gls3OZO
jSmEhOMP6cSqc75ulmNBMOcrIHCGlSN3rhpqwxK9yS3muiANg86iTaF0C5JvqhTMUrinnUTgkuO/
wgeSAI2IXR/COZNCXp8A3MIkOohe8gP3sCnfqsvQkebwKGFeYuPYFJ3gn6WxrVWJGll5BDyHfpOG
CFMKdx9G/03YtjKdNJzzugXlVGMxWWU20/iOp/j4aNqFit0NvUjMvTeK2av3DonwK1Qjd4RHX/ZO
yciiEESjQydOSlcEYNzyo7J2ke3/3nsNz62f2U9Daz67Yh/XRCBuPM6qXsJf8mMWNlVx+wHsEbMx
jiBhUfAzp48pCD3X/7QAIw57h6ydbI+04p4krdCrr8F/mjR8xMkkU++hcTBz1jXz0qBGSAyiv8oU
Oz5teQZHBO8jtSCQrFl/zw+wX4bxkBsO62Q8aK2WRVQOggzlnhgjVq5NES9bAE06y0g94Fr82F8G
zbpix7XDIkQZIl1tZ/DAEUc7RkfJ2ftP+CSx1biWOAV+EtYhC0J6FXnts9XrYXweSHDNmmRmih7K
dwBs4uRc61nCuHRLiRBWaxnbHCYTf7CCsOj1ivMHBVV8DFl0bwuB6qa3uemiuBd4G7eeJNsoEodL
rUQqk7rVToPNrS/Mx4El9iREFTMlD0y84/895yadu1gJ4OiTxhYxX/BFu0jhLt9PUG+/E/xTj6wK
JTINLoXRIq4weJejtHGXAsXJcTM6umgN0LrCPFzKb8jcVOX7OJsXjd9EyLEJCII1bCuSoeNRfhEN
FyCoy+IiIQX6s2ekDeVz4F7QaQ2nTNAOUuEtQnJxfIuZRo+nY5w021s2Nsxq3IABBDYiPAu6Eqn+
GLLhbpOIywcl80YhBI5FlmjddLOU0zcK65zEXgirPf3VPN93IT8/E3kkI+ALbsd7RmrpJZVO0HIo
UDcIMo34rk2+GD3tZWRspvk5AgC3bKq7oXLNOwgtWwSUxLVgdvaU4d1/hhm+aTDVK+2q/6d+jWpU
3NNKjs7bpfziPn4GnBPH6Y0BmSUEK5f1643qgDrCNI4AjIdfUFcKjso4ade0JKflSVwJZ4iANXEA
D2s2gagX5a2QxCVh4pIYhIl/vop2mM55tk/tJWQiDGXLbrfXkY9RtkUPiGuLY7IzTfgbtBOQSgSY
a3Mr74B4gcNxCNpc6Jf2/A928m1HiVNTWk4+jIKK7HNhl0WSk8SvzElqDcOxNX502Jt4Dr2kL8yk
o2DN8Eb/phmlaQ0v89bBxAAGuN8duLJMNEQnIymjzyjliefzSIGxSxRjlT1xdZET5CWLFIR7elQ8
DLG3Q7aWIrerSHuLNAC36KgSWedIRf+c4eArj37Our49K92uF1CEhWxlZuh9Mo6E+GLKGPNBKLJP
gxh8CqrpOqDf7prwTp2QdxPixo2a9KERs5YZPSXnzbamN+WILde2r4v/LFZQL7YnFxaaozMo2K/a
n2vyYhpEsi/ybPkqWyhJwlGoa/2Czble+rSunNArfRXSSGPbf/6tLMj0XUmfztdbiRUgUgkHAicF
Dbiidr/OZXAsCnL1QHcov2uri3zBz2bmXiA8ZcY4rq39E/z+CvdgAVZwtYhlztlEzWQUcUQTmLjO
mXucXXrF6/zpFP7lofsqa1uzHXvCa2mu4KJ2PborOUFnOhQiZ74UgT2d90sjVmfbaNrMODF2Z8s8
G6yQMmrxFsg7jX45/GCnsFSfFaKL9ULKTHIKq3hR1ap6BJ4k55pVKJkh4Al+iyZ+HU/LCQDWc4j8
6pNEs1cigkQlIbODNZPivErCUMluPF88guRdqpzSj6hgA1p/SajEZjC9tIVQD+MW6p8QK60w91UX
kbrT1jtoxARV5BlXhN42xhzjwQ5apOkL+NUt3a1KKGc4vp9RdhQ7XxDWw3WI88WmKs1dwIfdgi5P
U2PMQGvwt0FL8B8Y/s9EQfR++TFrHuhWrOP066/TX0iy8nqXXfzBO0yAot3Oe/d5zHP14rkMobYc
o9kPVlfYbWm9oUtUqM6R+0Q7YGNKBltEgGPQ5UHj5XbM7fjE23A8OCN/tbiISEMM1nE0nuAfE9nm
NTXGLoCHvhWSu1paqy8+VhoKxQZ4RG4L3qk3S6YzGo4Kei5gMod1lnRDsnHQsODxqPpXvBCRwemg
ainQpZ4iip9XnO+e41Y+CRsdcFaM6h2O6lDRN4PPERLIU/36vdrw3qHuBOcGUTaE6h+NubYf0JDP
2zKDmPHsez2CYkPh9djtB/ZRagMrouvnaQJYoYWo3RVzASg45TM4SrWA/L4P6gJ5dMUv+DT0AX7e
8TkI6jUpjGtAwTM+msLDKf4AQiXaUdAPWrDGG9M3NbpqSA91PS/QynEB9KJrtOnDl+VbLqA0eP77
FeKP2tldw1P7pZtLe92XclU8fRpfhByF6RDd41HXDsX2kavH5sDObdPEVPsFKqRUrkNT+3H3EMgG
wGloFHTVSxG1NUwdOr1U98eCo1+acT3Ef7pKDqaSw4mgZXbhYnu5S2q0xBNL+xp6q9+FGlHX5ipi
ny4DNZjYgKDajxooxiECydhLuIaCrhlb4HkkS0WIhcIErmosGP6imXBjZdKNIqHFawaCdzW0yfoA
MbaCSLplK/3EVtOCuzv+2RUXZZy0khi+27UqDeNA1yZ4FFe3yCHrqWHs1k0wJOMr4BHO7BWOGgaw
myoiCjPqsX5x4fGulrH/JJZCQf7LRG/eOaX4ogAB3MCW4SpD09wJPX15e5MxfW2p7dzLYgxIAmRo
g4emHCbLsBElGumSzZw2NNPy8MKv3/6Heko8JdaxlPCd7KByV2L1Oo1n0HE11E392qSDxgb8Hy1k
wrl4zNAmN47kAxfZF8GpNshPnlzu8dBsLX1Vlw1A+4gr/frhrrtszKjLI0DDHCuAR6Qwgg5bBoT3
fyYvlcgKtTf/Dc8GZJLDr+UBfGhjq36lzgKqQwPeEC+d4Dwp0TQhQO8UNUQa9F0CPFPSRum85qDR
4U1MG+3GbLEbG6TJHm/aSaK+fgjUv0XjZ9PPBb3A82lE/TWwGmFVGW+AAmCgIS1xrm0DXvGkEuZb
n+fV5WtflPGP9sDljJ/wdKnJ/y9IRl51oNwD/YQtX98C/NsmsHQI4Uu+bx7U41Emg6+/0sJoW2AB
rFPXfAyd8lBL5PWAivzs0AhRxlsjIodA1AcwDkCOo4Tq7g3V4D0QS6tZJZFgaOVSaVfrcSxIsKfe
K64lgR0MyFtkfTAaQHTJpSqtAMkGX+iCV1uKQm5G+b1NRp4VdqbRYVlojhAUoKx3UmdvAq7QrwQ9
9Dqh3hxkusA6RBWAVNgKoSfcNgTLYzPVJ4jjQQB8PFgl0aAObhpNACK/mTs/8t8YQBmBZ8WoS/Ey
GX1leBGDNXEFnRwbOGh3QHsbKWRWb9RM41jwIOQsn0ZyyUtVessDWdMaagrYRuJDqnv94UsEu9DG
iYcU0FdRN+Y+13bJgA1TeEH/h4XvGSqEFdKiSj/Hkdc0l5+q7/Ahcty9To/6AUQqsHIIdGd/NXzO
HgGQ6d9qd8N1dqBXnagxDfDyT11UrJf+/LqpZyHbxxJxLjL3jBCXdB10l7yTwSWtsAst90ZTr/KG
gpzEXFoPUOWhmrQKuxzic/1HPON53BNsztQAzJ+YLq8M0Uvis0jlTcWKxCgVtV3kuG+FZ/ShZL0h
Gq/xDDZOhfCKPYpmywsoAYRRb9UzVRI1AmUXCNI3tej9ovtLsAIBfjKFaZfIlE27AaGKXs+WRiTq
QA2JspYfDGOTp3xihTa2UJezbo+5zsCojpZCm6BgWrUZrOqzvgm4ceT6yoYo+QiPHIJKOviNksK8
PoAqp8zP5GR89A0Xqfrd3cYB3l8mbMNxhsXrdEFIkmzDmLVYdNIJlqbKwFN+75+Jvm3sjnjDdH7T
cCBfvIdhO3OGilZAJGKiSAYsyyPPl+jQYe+iJkNHeH2lqAnrOW0f1hlYG8Z2b91gZqkaV5VJuYDr
ee3ck9M+pKKs11gVR9Vj/Ho7Mv7D2UcqaBn2hHpV6sZZBNW7AgvPtXi+dCHv7gOhoOR6+OUUgebG
rr4cGcXHuMSgd2fZB7/s/rBus+TD04kqlXiT4XuWEArtAoQkCAyrQXUWglfSNIHJqXnfnjRYdl62
ZYSWsCg6t7+Zuy+E9SjFR4ld0YqDJBe1MIS9m0O3ac7LZG48L77/XIQNmQ00dijfqm57L8rUaP+b
EUnRCx6445EeBWb+KHX40CcvGVaID72CyCdSlnSMsiV/rqaA6JgdH79Jo50dr64akJNeN1sD5R/L
Pv8ITM0lniNIMF0SlxQDWiSalCPiLUJzI7RncS0QcQnMVlQRVoG4qPB3CQxutbcekM/N+FwWqmQH
D6FHSlF6C247wJHlmgr0I3yT+h6PrxDqClaDZY7Z5ZeZuyoKxFHSgskW4SVafown1ORF3hK84RRM
HHGoZccoW7Gsig/M3PMw6gjS+aQzBJE9oRXu5F+/1EO4Z8EleN5iPxXX5pBpo/BJCdbtXtXBd7Rd
eG4pORl3dI1/qNwll7uBhVwwHP2Bm0L37+JuNBpi5MEUYgHQU91u0r+zclWUD4sjBELtnGwWtFO2
CfPaGv75rHRDoCqJAXbje7eHc8kbg3Tj9L4n50GTkwA98qTgS9/BtB5V9ma4LrRiBsRUEcbpe9oN
6q5oAsW7aH/UiRM0GaQUbV5J9IhbVsYwQKr1rh7r3sHwVBo23Ra5JrQ6x0I+wwEmUqFYQuJ/Sbe/
9v2Qnlhzp0NI0TjmxfNJ+yKdCECmQHnfIBysqwBbbXtMxnbZH7lr+oeZAVQ1k16GKo30VlEuzQ7J
zeGKgnDuYf0RFPafUx6u3Bme1TmIvEK0dRmL3DAoV3yHVH/GU2ArKih31PpYnJjXknpgLTsEiXu6
daydJL9O//dphC6fOtixiGOWiWullyA5zPkVkT/lITROi9R9BwNcKiTe1nc9Zh5PSr1eq5Zt7g60
b5yXJGQtYiOwMPrKRQPe/RzKqHrorh2/TGsrLyJArgZln93uhW+vP2b1qit4ay0ubXsliH2CuyYX
uZnBpYHcnCLDGyrM+AOqKQEdlxRyR+B7dOCfKgZWFbiERIii1xr5UW7OKVnW8gSkyJTC5VVVqm90
xd97KQehj5PVTZ0ph/6Idz29Ogqntn+WABXNIbemGZ+99X2t8LOsIsHZxa00k3lIz5WZZACWC8T7
kOFB3IlLHMPTkrXu3uAcXdlpvGdK7euwcmw7eujOWicf+UZ6VFWAOI0MqPN3Jg7CX7WZhubms1/N
1tSrI072N1M0oDxZt+TCyLXKPLzCaljty8T5mY0xnZPp8oWF9Ppn1G7E4wI3CCMDpBtRTYPPE2Gc
lfvUDq6BgrQi2ZQV5hAz9zpVSDTESN48gK5iz+uaongHadkLKOAGvBMvunBABPwBqhdl52Hjt6JL
qD+Ii0wfG9qCHQB7RIkMetF4nipabOwrFzlNH97f9Uimz38QUiq3fV2s7tsKi0R2g+5fwqt+nt3m
/TaqD1/+chX7JKMuK/D8KiL2ldLyq/WKcBaAHxtQfuy2EfG9mUdTuifRBLCO6Cs5Vau16fzqhItn
9jsAnsvqMZHwhufDlGa0jG5G+aZUGX5vdcYeOFiEoSw6QrGuYSkcTWWOSFZPNjoMeAnnA009uqI+
talrkZj6yPO4DDS/UIMV61LZTu53rm5h58PSh7PB3/ywu1raYoaeLTlaCuK4BS8RZ9dq7stfAPIp
rydkVHHy3cR4Vo77S58DEbW5Lcjb+HqEITkDMkHe0DjKaPQwkj4F9mdHOm3ZzCjX+BTuZv/kyNtu
DfY4eLWABEmYodzzvWwAPzSjNukiTeudilQngrS51obkLKNnWdWbkwpSZ+wZHEXF/nAX18zglY2k
4xoD2enltycwxpTZdI8SnqkiBQD8v2lG4obC3XUaqDd2WV7IXGXRgv1d5Nuf8q9wolCxVCNTMwRD
lPlApxGCCCxSjCb9lRR9vG/ac7lcLteoMAzl/r2rSnEfLN3u206MFVXp1HGKAWGFvYnN2Bnn48jP
7S2cyFB9mQc3ignnSjr1GF8txNxA3dfOrdFeqr9wUgqj5Ws9J2QYh7Fe0+/BLtD4vNN72gfBp159
SkTWVK/PamNGC4BisvmwFKtUVW6Lk/ia3fMjfnvT57Wqo6Hq5i0lWx50pgJeUoXI4tE3VKam9TKD
b5ZIup6y8Htc7aXc5DbHVsPxha/keTRgdzfLqFcWEILVGqzIeYVvtCDotAgjp1A5y2miOrwlAZN6
Dh/69A6TsjFb8MRDPafWgEZBCJarrW5pi1Ke1xEwVkvd2uuT5zGEpWp/YTDy+g3fkcMQDFpEvVws
hH2J9rcIdO7oQWoqsJ/weQ4irk25xDklVsNVXpJ6NtNZ+D9EqpYrZaSINla8C7b6lntovTG1Of7J
/TI8yvdHOqO0NuiNm4/7NgX9zZDvlvs0dGvS+L5aA0NCnz5jYkMrzXTRIPzngLZVQwulWAUpZP6Z
WWc1NoMNkiVE2R7+mledoZz+1rPorJ3r8T+f5jLT6EtZjvojiT7ZnzYGtXB2RIx1Wsqb09vewJzD
q7JDuVg8+3Y75qeOfr4kqK4WSbSNn6P2pCF5OmrtiBR4nlOWNDLOIabeqnlskeeMHGJc365hEC6w
im70XBLY0LKwJxS2PXSFCjxXRy0cFvtW6UM0Xh7oOZ1t/Fj3GoqcUnu3aQBgc+k1gr6SZBu0udxZ
qTXBHZDkaUcCrO/uoipQQOIieCR6+hOanoxYBYg9/3/Inv2qUPS3dKFveoaling75gpTqBY/b/WH
h5mIfMERJ48bhBmxdvDxZ0bRMZr9xRczwDZmDx+k1N/IOtoFTzuFLMdduvPiSphn2BYfDojFsO4P
pp9YZOOGJOzG8aVQqvvTUj8evZz0Dl6Ocwi+Vq7CKUX0IeXUKJmOO0tOpEbdfTEbjiGi2JvA6zZ2
DAkE8neoQXKA8hEY4qQXRRZDBrFmTlRNezfhN6MqWe7DY60CatWQ/sqUY0jg1M4TUobTRSDf69c7
2SnX5AAhRKPjjzS/erDkvD3SN50foQBgOBoHzVLEIM9Yl5Pugi9/8VncwfNF+SHTGbxccKVza6Dv
dpY3jQzryOIFt6/o4O+ZX2D6xTdbNVNLSjXEEp3galzyI+yYb4rSoCq3+GaxcbTPoQtRhJgubopJ
rQQ2z7ST4Fz+pIUAbbRM6no1WFV5qiJEbE79LFOYXTTUYNMTtbAqW5cjVKpjckFEE9BKZKMOPbfj
8lejS/QFQtDyj95ABuKqpn3wKxfIuFBhPee8piScZw6wvMjXDdL/NyoX5GoWEHn8t4VNJlzIzMFJ
WdIbOsBsopfvjkxUevzGuF0tI9dfbVRYK+2bS2NBwyaKZWitF5pEObCDjpzUlC0+1sKQsJwx4phV
umG7i/IM60cd13MweLth1SbL/RI6TyUdR5HWs6XjfECDSYbH9Tba6xtXnArrgEGvbfxkZ84cY05R
Ojon8abqW4ddgwb6VoPnZX8dGDfE82/OdFhYEq2PkzlZcXSga6ffmF3s/h2XH2VH+gIY/xYw/djJ
KM+h1ASr4wCrs2sqj4hb7ougRUjRORas/SfLxOQxDYWPapdQg0MBLbnVl9TKXY0iMPvHwdKXF21i
f/PNXL5QS0b91d6e64AOrBAKGm3fvl5o+z3A/HS3K8RhIO0Ix2iL7w6oOz8Aj8yIWuFON9RfaFyH
uMzIrCxc23iNJKmPGvfyCZzS45Zb05/nzonQYiDwhe2Bq/GSHc/JZuwryMG1hwwIw4KPwGcFIGt8
ouoldAgeGxbdz6tawD4Mu+KuGxDOAv22MBadm0CgbuJ3TpaTN35ebvL8nqE8aI+u+Anc8ADa6WnF
QIx3J0/yQeQ+RX8PfSVUltWqBDT8fKZ2D1NJgkq/ws4HBF9kk39h0peeuixVALYXT5GffTOoSEx5
C2CvhSJlcddT3SKmGyrK8fcjxEOwOC4MfK0mOz/AYsnwCGtX31db3ECRlqt29P7U/85jh1eoUH0d
5YPLRth51/etTc4beZ60NjrUbV9GSWPJ623y8PO6+433M395C9PPOVZ9/BBt5qwR59uuqUpxZlXt
181eIXhJ2ivK1WMBzg5G/FyltuDGMEFRNULtbuw60+21QY+/RkrIDBpZ3Q9wFSogVkraEbkiGHqm
/lAVgfARYfbSvJqmi85nYgY43tCB3PxHB6I9qJTUTAteETApEEGKcK+sfv8hF13buB8m7g5LApWC
JHO4K2Bz8+ZDO9PEAXCfNs7C/13z2gboMU5cmOkMrFb8GyWO7f38BLK/X4+MCNHdFvp79/kOgf+O
PCTrKzM359IEMozIZSQYDIYCOdygjP/zhKnVQpz8FeJH/u3ru/ct1/K+sNJtqG0yyfR0y0EQLt98
V1NkX8Nuwn2l8XdIXuteGh8sD7BArw5u/+GfhJkbmfo3K2oEmKCk7yN8ztGKgRNaSOI0x+2B4RZE
OFZzABz6y6PbovsZNQdFlzsaa86ab8Ehq7p2JmwvBR3Cu1yP1v+A/jxXB3jo0YjERy031cJY1ART
ictLhnb/hEvKWtUbextVdNXzJCADxHFJtDljlFrqzkRsdVIi3UAWetP2gT3JSDVynAeE3tf+0Diy
xpcf/N3Uai5yXGyilUtqDLxwU3WXOF3d8Ue6EO3xnfgnVFN4OSDi2w3GJS5a668vd343bVpSVCQx
ki4kcilW0+pjwDo0AnFaxoy8SZVmXh43pdmykgJLtTljBUTDRpwJ5fmVVOv4kRuZBX+W3Wim72rx
FJGsIR2Dzk0LXQKAXJmWUloobL9+53aSdAb8EtY7wRKdmbhmy6pFvNuxlfVmASMZnodQxgN88N1H
VJRHSW3lefgNJj++aM8tIsmJu9G4BXZ4Jc5FNyvBW/+CCMBYWLWevUJs9LX82iKgyXaKLUf03lbi
tX7C7obmdQ97j1sJKwyEOzPSjd7nCn4y1gJH08uxkwuW6rv/6g7uP9tF9BLRBXuZ/pIB1GnaNs5R
aJXaTFlBY6M9TdHKQLzQiYywZgcj1SPDwAP/yBAnjjufchRwYdlz6fwN9lrv6RL702DTq6S2RjK8
mYQtcDE1fC3g6DAAyfL0Ega6EZbxFuVTISmvOoYVqoOEAXEdrLU408x2PQjzse3B7z6Ovz244e/P
6mlYWyvwAY2JayPh126J/GRfDxOaimDmuWNJb+2jwhb/1lQkXDI8nvOzmlh41Gza9/UEDPFjiSgi
SUdRQ2xO00/prMXJtB7WWrT8UBkvtAw9GjFkitfEUZl2M27FJU0K12wRsiNDCa6M9Vweq6g0Ei56
8kmaSxEq3DFZS8FvHCWyKJuOnvrl+zJ6AeEiHGzKGAGVyAvedOQo8NBgPyDDNGBb3KLUDJcbx0T9
NgnbbZiWujfRdQfUTMzCVcbPqWUWC4DDThsQX/KRgmCO8A794KOjJ0e1TDUwLlybZyYk8yGYWiQj
vPM2GLnQx5WVErk1ac5ICwgCACKfxriXncDcs65J+mm6uO8mdjKF4kn+I5dhdRUzJBOeFbe3pZRv
TpJXPdD4yt1vDzZT+CGZdnEof6VMETb0WL9hRFACC9HYJjaR/tDU1ue5ZJECeHD1Pbp11CHXIyk9
/feBUCIYcG7WI3kBF/Y4GzO+KDHwUx26phhfpn9eymyQmZt/JzOssHJiqRVa/q0NsU/o2p3/xAbd
HL9/8S1hLLu7HroOsb9VvNQhiS7DZOEsRTY9F+Af0dYfpOMZfANsFhD1VLZJMELyP4L4NNLWQDSq
wz6fFq4Lj0DcYkflLIufdk3ags7Xetv3VecKPxELJ/072+zOU6vN0fFK2ZJ4j09+UxuvWyWwIlyt
RWKi90WJQM9V338W8GkrNzcHWz9nIEDs29vyWEVNk70/8JbCqwq5z0pH2cPoM/9sZX8SQI54uAkb
GNlegshYc4Udtz8p6BsAu+RMfwjHLCk2tFq4PqWhsNahKVBAQrnDADn82veFpW9JDpA+5OgntNDD
wvdgB3geXFo5coBL50CUSdXdSZNi/gCdRWkpo8Xrm0QSvGE94qfUc8Vd1sFZU7oTkyqqmD69FRmu
5qeu57PsPT4o+E3wdWaf4cU9OdThbL32f7XEKeqF2v71SYqbsoKMvSNoUZWazduX2HbP5fsZGR1S
GJZhm4gi1IB5+gSS9ILH7GQUSE+jBCW1EzYvqyt7xpFwYhZxfzFLoQVsmecE+GYHDw5Wk0gpfPaL
lsaZpG7UfeiLQlxRmh+3oB+zK1P9vy/sjcyu9HPx/Wahq1SSGRaqc6RvZWzbMLOJznzFsNnMosg=
`pragma protect end_protected
