`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
OAstTLBlkJxExOmbDz5Bl9uqf6jyx4d+ZlQZ+/3CnG/ZMotM8ImmEL7OhF7xffWl7pSBwds++VnA
P3tw+ox+XQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jx9bn0/3gtr8IYHsY3HyDX2LX8tf8Kr9qr3/pvWBThcEcshB6L8F1LCJMOp/h0znHOb7DI1lkc1f
fpSQms9kcrqL1uQPDQHIxamAR7FkyXkOE5Dtvby3jtVIpVf2t5GlBHf+ZMqL+RMzU6DstDC/qp0L
/2/n3Zs3QW1Qq2kO+Hk=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
rZ6Tq+OwGsTKXg0+c5SGURPRk930c9FFjcBT3Zl6HxTiPjDH3U376EVRKm3LkdTSYdtZ0Qq9pfUl
bVTq3sQ4HRxNqq2izWcL3Lc5qAdR5pE3VpKsS0dNNTkrsyqKq1D0/jPpHtd57deyom31Q7N2sMLz
T2ObMCNcsCRQBbgcaFw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
BhMbd5yJ67eQrGpGuxRO05lgxlxUcsmm1H79RSnqLVDHfINifIcPcwTh7rQ0BYSEomlGE2f4xjTf
Mfz07yuATc7hViMAkCX2sy4B71pQHOk9UVlgt5O9k3d7iV3BPl3CXYg9SrIyt0ImDFaP7uJhgXQK
/j6sIgAQnVAmr9yqpvsB9s/ARi3gP66Z5FOf79TX5o41YrTPticAzfAdDv//mI/12PDfiFucWHCE
85b015PEyQlE21+hJZyoDLOohNInFecyDy41h2er0/tCpxhCt5BCvxNgVAg5/cbl6apFm6/QTDms
6XUucYA3p16J8OtYs4INeLAk2Zt/sl/LkIrwnw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
F6GGFG2GuG1Tv8QeZKiJDjR7+T9fKlCIAEvwEmqtdO2LAkheAhcbqrBi6RmYZKzg8sZBbIxGBqwy
uwXr3WD9EYcgMXL7E1EwMMi2CgXkB0xJjwUbkbQiZfJxaMKq8BDhJLwU/PmYqwo7fddV0JmA80bb
yjpTTRptL1Jpqf87TRLaQ0ZmtM9kGMXwrb75YzUQbAJnqYs+Rsi8DmXK8xbZQ2fF4E959s0spckX
6uQm4ACVPYVstbjJarAJ29aA0d32Cix/cf7/5lB27b6h8u93oSCGAB3eNbVUBsbj9b4U+d4XY1j5
nOeJmchyldRbnMHXMxq+8OtajAG0JrAN5WFqwA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
UKtagqMDYxO/rBPiNirWiR12U4FJmcezp/KPrXLnn4cOYz+25bArSvUnqomk46HZk8qlvhkDODHi
EZ9bj3BZ6lYlUZNT1d785o2kVu4ynLPaq2EcZ6sAIFpq7RsoiGxJvBbXA+ORuSPY1z3sdMQsfVMC
j18Z9wCsUdSZn4sT8qJx9i/Y/pAoVyNQTgGR2drylOOXIbHcMIkpDXWU/AtMQ1RBIHhZyvrAYRRM
PQN51pqb4dCj2cJ2JHFWXkTPYzKCYewS5Kajxh/6e5uTVGzgfziYAeo+A6RAZhYm1s/2B6u5ho43
5VnSbtZwsDHmVRPwuzB7mT33DWCiOpprnqyMOQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 151824)
`pragma protect data_block
7DPXtSjiC1xg6C4hg6hy4v/De2Z+1V6GT9ENWSO7+q3fzWTQgI1mULqlNsxao2ealg73ri+kWQJy
9E6tcsHr1CkI9kxCD+ITgg6v8+sHAw8TgD7uJaYoiEWr9IoIVKvWjNVgBoLwNNxbNx01ysUAU9kM
jkUTdnTr3/bjB6Mld1ZMaZdIExENKHcNKwA3I6ECKc8+jcQ1y+bPDjW+MIB1qc6lL1ep7J/wb1g8
rRTTH8+iR7W+tyZl+vG0EIcSbaeAGKnBQF2XdRRtOlJODpklBqE6tS2QUjZ8OBMcspy/vKBtZyVR
J67mOKUir7ip8pCDVfqLD2cQtMGF21+x+qp4GoypwUhHAMi4sQUw5F/WMwgjHiDhKKSsHgEVX1Rl
DtD+idaPpX934g9mkdR0SWMX5PG7L45c11kCZcDlEuAG5u/QlPEQUJu3WfS26TZwdwIwez5hEr8J
vtg7Bpakno4/z/b7hoEdicwqXo1tjqNJ8qdC2z480zT6AVhz8CrU30DuzPR+oyo2K/R5GhJwkTD3
NLUDjJzgJq8CGdeYSxHe7EW3lTLKI2uNHM8nzKAOWzurYKs8FE32e/0eDBcHLDiCb8ZmkQjnSxje
g3rcgF44s1Sg06vd/HJEec+jvoVP+hWiJl6K67ycMofrxGU7pm6ajoxVZUpitVBdpd1FUwKaC/uc
l0QmMhItcVitN0UNHEvPsI71ngBPjc05z5ztnoB5cCmnMdRwiXjP3sL0hNFoX10LatIUNvrvh8rb
I1MVtSmvc9JvHm+zkAstaShgnTwGtVyptSk5Lp27MviYhkAYanO4nfI8O1xzhYJj3dPLbeXsq/OM
2tttX5h3wcP/RNlGsuVgVOGijrlbMvxKsBU4CFavGPrH+DEiqOda08IEBttS93ANIlQ/UHIdyfry
nfhKlxVYp/frys5lOCNnT99h08cpou4e2f6IGcl70PjQt90eRKSZM2AVIqPc3GmGaTt6oQbPvvIu
dNKPG4csyLU4mh8GyucdKyOkXbrMh8nmqCbshAaAc05YPDSANxBX9h2nDg643ZxLVDl1ybhi83yH
N27i7VQkQiVBBP9fQPqti7Apu8k+GN+wx6+ka8e5k35WIVcsrlcPxJRTURAI8Q3sh7NSB9JAxs1h
SD1rm1hrEk82meemDHYt4VxxrVBCFUdpcq9y13uvZ4XG9c/MhghAoroodhiQuCqUH4puGAUXKuoe
n7YUrSsGwK4hpe3hqAzCw89PQSPRmVdyA9DsAwD72ZzgMFmHvKHc9GWU9HdHjIxNAR+Hjf7kl8s7
GggPzV2da0u+D4Q9XVqNiiURzvwHPXV4ExkgadXxQRPS91Sgw9UCSXyGUz8h76/BqVjr0rhW2OvS
tOv3veCvsCHhYARIWQMP88r26xDNMm30g01oR24cr0FDalHN62GyiMN1Rvaso+1ZB5zFAXQW79LW
l5wq5046LoC/Z5e/39lAYCkJcohwFoM6SBmCFTD4Tb2dowun4oMnmwG+z23UA66wnE0VUjZY0QQB
WqSQy4J8sIAam/UcIPh//kSQC3Y+1iWWi8wVTt/mH9RT6QyHkz948p3ycQq8XaD/LwHpqLRimDNB
Icprz/Zvf4lO1S4NYD+1gZuxDo8c+zzitplYvyXjE8wBEVYaqx+YRWkirNtHjgWVX/JmpxBiNUtH
ywPTwTleImubjQSQOcHVC9sJ2Ihvh28vN42cvqYPcUtC20dq+NOaNgnQrjNUXOJvAs5mMjQjV4Uj
+k/Xj+dM2gNTSyRt1TGCcDR3rQMdF0Ks4d0IP7N0WWDBB8FrX24WQSET9oh/sQW2RArkstkxzYqL
7+4fz1LXop+RysromeK0d6GIzUHw0xCox5/jJWH6ZQNx0ERc9BIjLZTILkf/62cA3a555iQVR62j
BDX+lpUg0DBE4VlJjO/D7qwQBOVLAoCflf9V50dpH0Rd1AL72657qt7rtMLrNAVNdcfZXsdlmLFK
hU0sMs5z5zze7qkA+D+ZM0Syq3scBPMlSAJLzCjcGNGUpBuobwGl26ACvJgZZLaoUXB8eGzPBG3j
AyVMU3S3ANuAckFXoSroQwk0H17PXRdfuLPb0Fx3gZSc6YfJdw6eAiVgQWH1yNswB8pipttjrg/n
PfvEPDDX98+Dv/fX0bQHxl2fIbD7lImuGn7WAu8ClpFJxPPBWqlyzozmGx2uywcyztktDPCfG+/R
liomCi1LmWv62xaa3AWgWIHvSgzXW+JlnhSxc8jOiGZmUUG+5AvGRZc72nPXTThJUfGC9h4eejiV
Ho+fg18rJxdhziRoePXXEe1FM8i0sMKS5/iaU4SNcAB7JdoNJ+0E2K4DoEGDcqOZRKt4oUMtuDUn
IGJYvvmvFd+QdTFbxNqqHci9wVxwK7jKhJZ3eChFxhzkfes+hd1WJASiOCAZE1nEPlmIrUj+jBm7
9cbg2/vfTdZ9LQ2TFhLy0ZazxkS6drG4yKXFxYCncb0Lu5agTtC4bh8BQExiObB8TPPsTzixhiFJ
c4HlMuNSjzzDKoV51wjtvPq5Qsxj/ylgJJZvn4egaAKcc+vVT0JC5eQjM/3HtOeiSPcgMTrXkWy5
Sn3cJB7eGAZTf1Ac1aTvoKMq6PMKiIPbTQwLo0HFgutSUK0dHJNcMEjYopJ5QJV7uMmjxo74qclb
kWflEKAFKUhoi3a8XOiRPObGVvOZTvk9gyeiSacvv2TvLxz2Vv2tIQA/36oTxB1VX/zUpBr31wKG
zSPtn7j8Md8UNAFMOQVHZEaXVHFgRK9C5PW04m2wW1o9/N4tzz3AJ3jxBUZjOKbQ+HrB6y8isb9y
G5cOqSDzWag8mCLnCLsh9ZZsESCtXreEL5/hVUxcHCyKtb7w+qX9omA1n2p6vVQ2M6jwJX+cLjie
/8jnG5PtQllhN8AO2a6d/GbGqxiyxHi+RE/F9vHPUQnmaRkqUtVG4UUWT4Uk+STR2IPXMbAO8W8o
iIQTidbjhBPrXmeO23VRys2Mu3QDjFYQIGIHsZCLsWYaBJ5d4jqev1aT24e9MerAGSbCcE+/mVyV
jZupxkK1QYbCZylrhnAMuUeVejcw/fMQuza9UQ3M2lz4y+gJcda2eyDjmgG+iHAroIgywTqzDDDg
csX7sqwdx9lVZvdGQNVeAAqnP2hvIZ5DDWIW7qa/e8SJc9RgJRvEjlgaAUM5/jC2B55J4ZgAKgWb
c30cjIlLesnjKvOnFIsuOi33FbuqoP3MpYTxUm88VkqlxLPMW2SObuakHJM7yf1QQFHOxR42kwa5
bR5Wdep12gcyboWxtbPF3hWH9q/3ZnMLeXrcfG6kFg5wd/7yTdVMH/KCihA95EnEjNw6xCYNuYuV
eMhGZhC/MdGSMMcOVMyY/nmbhkkMTVb79ZNhBmTvri9wr3akdTRKMAriJ4L1bZg75QsSVzaZ7rpQ
Sr2eZSEzV0nAxXIAH6DuL5oDVd0iXMA/gpZ8mVz+EP7S6GC02bi2J0po7hm9gWQ0lpSiCMGexXjX
+HaO0IbFV+K6kiSyHr/UvJITDgkieWmDht2ccRLok07VR+MADvJghrPR0VpOWZB1JnNdJuuR2WW0
rxFTJjVF/TZHWFjbzgsWMQ+UdFsJyrq5vkxGhpnk6NEtflWNQvPx6R/Tl2/ZNjbg1KT/27KTDgdK
oMZwtinjJnUrUqkVvTvmnUpVYhGSoViEwf6Mjj+XVTlN2WpNfgTpS7g9F7tnpzSd4xVeXzuIMnCj
ExObMnmJEEQvTs+ELkW+K45LlBn7HFo/Pxi7MKnig0FRYYBB9hdAJQUZsXafE8rI0geIjd3b9I8d
c3zfFwNLcJPwFRdBPNUAy7PAisCk4XML2fFIrfe9sbH9em2JPHftw9ebxfVV8s5W+IpZRYRqD+WM
v5wWaNf36Pyx+kQHKTZrO7dVrDyzKhPIzamKn0vWgDfKOl37lSXshjXLZoi1qGM8aj+GYNdTAzuz
pz4e7mPgAwhTacBnKOFQDBZvwJtG9m3DTpoLrfTaNAJU/Acu0hEk4twQTHJ91ysGVtDyuVC7YR+4
od8aE20zEIomIM1AuiU5v5rHV9n+eJLteVtPebWYYFKu3/Pm2iiDu0EJKdvuAtIopVl57gjf7wVe
KRqO6T4AayER57Y0W7YXMvCXkOtvid3ZVvUqyvGFHS/XeAgMVEsfk3LIqp0UAR0FJsmEwOuFM2hy
4SrXN02JY1EmjPl9UJGM9drl8qYFKPEV37KaH1n9J7U2nBs8WlyCJni+W5k02ZZwFc5LGSvbtwi1
ua/1o+nj9mEoKBsP3vd/QoA39zGuG2qU/WXdlpsm6dKKxTM6xoDIIjv2kvjQEh91nQywjuV57Kto
/6iRp1FTvJBBSHMWVQkltVzja4oAHd5ES8N/qfyaXMK8MbQOfhUf003BAGigmmISEQMbBthxKUjt
WLOYHK1l77sEjF9H3rpf9KEejJZ1RKvpulPXVlEZ2ETNRgi3JAU4tfYu3xbO8Um+F0u+SQjGJdSu
Q2CZJpoh96U4L8lIZoIWM24JulMgKaZ6r0jhEcnkWZUFVbDRkVlKM8i/mfMQG0ViR8W7v8BaF6Tt
Vp0lyMxTDQjmJRdVjnslc13yvwrZBa34mDSzCmN5B8DLcwaAcsR/mTbwgrmH31P9LI80vngeCuzV
HCqmKPGWDABiq55eNI0IQwf3oKblo6WmzccrJTF/nvjlESAiTruqMYrZvq8eVuqtLDljv98U1RV9
V/IsQWu7CyzYoiS38qrLKdg0aHJBb+cNRpWMg9rPHFVlObuT28cnb04NSpqL1PJCUntu/2wTF6sG
2pz1e4bprZZmg/yJHUsPU3sS66Ehj3jdrzDGcGSAqWuSREss8x6xf15jbNPRnJ0aQNphnUydpLr4
49ReRCCUMJts/PAmtBeeqYbe+mHb95qBrJm/k/2Hz1OyeDQxsGzYeeWI/pMEY3/H3jVSV3CCWVCh
hHzyNrSOAfNJA3Jfx6jdPhX5mWj4aEk1YQZSCUQhUBy5w8AdDWBYATzPkF3IZuhOerZxTsn0MdCQ
goTONu/0jMDdGiUHWkv+GlDE2FIhrag6vPAp0aLR/dracelkXCyn2FuZi2Y1Ve9e4jgfhNxQTuZO
ezZ+iye0eVdPokwyA3WLodIr+OwJAZNWz/LUNazntBQyLJ9xrOzFjVbatTY6i7QniC2vCmJjyOih
ibm9g65zUlrNpQsNQ06V7+WE9NpfI8adDMWa2jBM7pRRIVc3adQHBgZJ5yo7nqOlAg7nBrQHSiY/
skhnpzqiDPKrTT+vFHxKHQ8Jais08FmsL+oub4cSmj/g9hf7sq44x/4o0y8EPSEmGpPeRJelr82d
atRMGz4WuQcia6p4Kx6/Krdgd7LCe1fkLJ7DOEu25Mw+jMsBTp4Nb8GQzQp8b+Xbur8HJVHNViJA
UYhH4Lu0p0JABoc/aDkJOaSBBt046FRAGflmRY7H5t0ARbDq6J5VHh8kwkJSIqy33MAjBwlpnqyK
7YahIv9fVG4GhpN4vY1QaNTOLj+mFA5OIWBVcEys55adxFewsU3bgq0mdJnXJLPlz5EjwCqhFlHW
AznSpSj55waFAqyvJQ04IStBGxy999GqMwO1Bwsc6+H+BbHXM5UNPdtXW7f9jz97s07IZAQ1R19Y
BZZhWzm0iIb6ObYCjW9gmGRJ8HJXYjoPuqwqluMS6KGn1IZyPEpK1uS8YzqcIRZtBGk7CzTA2s62
lTo3grfochZpanFZG9RQlfWV+dK2qLjJqHn+d0gLbvoiJTgUAM7g6+v0aUFyFbqWGNaFZskW3wB+
ph8g50wGFDqABaQ9QnKJFHc1ORlZV3elCgDT+scC4co7wQX10q5S7SBKxkke34+tNar4BIagJwEs
CLef5h7QzXx3GdaJJrgePcumKpbEhnOxLmMyk7U0Xqf5of9rzmyjQ4XyFUE5udmsfp7DSKRl8Cms
1l7s0rI5Tota11/c3mWTkmD32Amel1pJPnsQTvJmw6LS9G6ObyB41ZDDOaomvgZpgDwiVHOp4CL2
JhaoGNUnJKQJ7Zqfi/DhKGeX1smSQFP8k/dpHjqECabiOH5CD7XOsz/BO60Fi4283t66i0fYaVvA
tERhaQQUjHHHBxwG7d9Uy4Blfo4HwofjN5Rz06d+sCthCUKWdJPM3y2F/+Zf7FRyDBKLNkBSgJdJ
HwZi/Vmmifm3FxsOX+cEPzPzlg4NtLDxVhBmKyQh5ZIz6LtqLv2bmQsgr1CBqZ1HzU0KJCLw6z2I
NhQKahIfTokJ/Bvvj0194aex3zK5erMk+FsJCPdwhCtExp7uvv04Bf4ZDRI5nwnDSiUFl6hdiQHl
G/7MKCraEbYw7myXo6Wf8cYcnt8m8hTz69dWGRwcGS/Je0iX5F8hxwltS0gUaw2EytMbCS5vdhRK
iUOSUls7ZcRaQf0hFi6cem06z46c/vOAHHp9uI2QAv5HfLTj4O7Mj8W/bQwC9QMHu36PSHhaxvMJ
ai2R5Qhl+ebJfYfXxcYlZ0GR4VMB/NmGXwFPDLKzsr3MnljFb51+Fjp2RutXnw2vbdkt8HfmRZqN
W1OJGkMTzGSRFWeP07SMlq/JjwtHSyvKAHqDqVoRIT7rpVZAcYlvbzrOVE+n3KG6BzFFzz4Gb0/t
nT33sgj9oiOnoJ8xA/N4K0eKhVJv5FnucIXt/d1Kg5JYcfP0V4Y2J9AOotOMPnvBgOmCKkv60mfP
frGd2Xx9Kmhv+L5FPIvum6UiJu+Vs1HAJUcLYJlfUsmc1o4KK/DYQvyOl6RHgPAcY+n1a+hcvqsM
GAkHi3Yts9sYr0Xp5H0V5W89NzMWh3xDy31Rjwf3ql/FJtsCuDkd1KC4/6U4C+uqGd7MAsQB6A7h
KYx5GaaFYAcWrE9oRpDBnMoFCqVH9J8KylxrV6XlVQP8yJQL/iLlVnRLXbIjr2U0f0FE2a1d4VOJ
S6MfK/Qp/PQq4009mjK6AXIuW12v2BqlHBwWqMc8s0OSgba6l8ATbFqhbjv/zzwTJCt/7Mo/52in
LmXCBu+ooR5cZWXyKulomubiQmPEdHlgrUJjMD+B2IMlbWmG3LehwDQwQaPgF2BZ/K0PAoguHMLb
H645LJhqRg112g4/7NvhABKb73Eq7w8k+w605fpGm5yBzvebpLiifa16JtBNGTrIOTSiLvjwuvbV
dDzLOQP+Ois0YDvbD+OacR0w4YlJ8OO1EXBdoDvaWTmhtaXXYWfdhyHCtjLYmm0U2XUBClTRBqXF
mHF/uSjTas575D0/7Wzc11Q4WGAkAAD+cAUd4tUdmvQi3KqbKTtTDSL6ByygPowffVgUJ3dgUaTZ
920x/BIWyRIopgqjZ+CQ1is32rviNEU9147+LRBrPt4pMU3F4aGBSSEpzV20Q73XrsPlrW+T1ob+
q9dfG2rnd5TTeh52sbRi98VHGXuzZ1S095aJRDVW+9iOQ5gMjXyW5iOOQvEsK1KGhJSrh+r97URJ
edbjI6662uqcSCR7iwWYxZle1XiGE1oRwH8qys2I8cKaHVKvkN49gviK1adhrfFGy0KqaYMW0x5/
AJpxvPI2IfeUIGGREoJjdu6hJBF2K1S7/8ay12CNHAi8kVa5VqjYlvji17NiSWy4uGuT4MDTxgPT
1Lo+j4IvuWyXKYjZ2C3fN7G1ckYx1BNNKdU0qS0+pYLEND/UZxDu2I1odY7uevcxkqu6Dm68lJr1
WIgSIgiW57qQdTjgo0y/VmuZd3iVAZikJuyJY1SBTMRRupB/5pLGPx3uA0qffH3F2ntJLvyH84gW
BDjK4jIE9RI5np1Rk3jSYovxhaZb/DXCMRsD1sY8bGjWSf+rYSZ/zi/Bw3cThQwsi/RRsAwjOtSb
5WX8USkrCxWFr7qidzbUE8HH87z/YlKIR/TyK0eqA1mKEUn3hcp0ypDLDhZgk43CwNjVFvFx6OS5
enmI1igoFTpJGkrNAfw8kjUBJknmkCvRSuDHgspi+LpXFDCqJ1SZre2eGUNc2SEIPfjH4ZQtu1g5
d1vmkxokcKe14KObPHyGCrXe2FC/+v2EQwoo2fzSCOmDvebj3fSaqhP7ucONC1ClqM07H3GhADmA
0yaHTAGgrvjo6/BtwZ//m7lUvrBdo9lkmSxWmuJLXZHxHW9EQMFSO3DJH4fcGXlQBGp4ic/5G9B3
M7jpnzpy+bM1689fBFGuYdRKnCedtJfLSy8o8oZo7+z7gY9lIzFXYJIOdin/cR/L8U/Ca8VLF10d
z+eTfUdEbaQauPxJvRCzXlPHEa+rDspgxOXZX36UK647nfLG9jiOCDLFc4CghCz1Z63nbuurhQ3y
heBFH1fh9FERKIjC9W6/OifGHQNQRPJvXl59aOBJolfstpwa1qmBu/pvQts2Gv0kllTOnZAIDal0
h7pY76YnbLc9SnT2Uad4hs0WB+npibS2URQsJS/1HpoftDnOWlxTNZbG8lashbrcOEbe8p227Ugb
fv6gFEoTllKCQKtmcNkmhAguhcNvQRnuB2e6edfE9vEu/FYXZ1NQfHVmsjK26yKxNtvuvAtUY8e6
yo3d+FcrJBFMvQyvg/gPZzFMaJcxOiFSgcb5s7cvlRHaTb5Gx+38DTCipTtUXIAmHdDO/Ms2wjWG
Ct2GvwyC1SBALObDbuvPJgaxkfEFsSgPm3Jkfp3/ZWSGLeYEtWW910OWDn3PW+jwjDjz0xMY+kmz
30tpOQPTHIzh13jBSC3No0WE/tYYtYmhe6NDzdSONT6f3uEp3DxEipJRYH3D2xG3DI307Au/KSiS
C426wN5zVm2AUzk27UELwEqZD+0xtAWIHSqUCgz2hfIER5dE41B52y7C8FxpQryq6NT6NutuPGrO
MBWWKoHxSZiTOhCGjReGA3hoyy7+/5Fb1+zkEW/sEC4ZVZwvsvFzXZMbsoQF+BZktXAX269gU/82
jNSoYVuT78IYSfd6ticz8nd4xojuXqW121x3bKsc3hjVCJOrO7Sr9/8+Fjp1rWOPaFxstImZ4uLz
atZSMaz2ZbUNGfM5y/RuDT7PJVrYK146rVcJ/PUAHcbtPUGx+4/b5KHCrNK1mm0U9PDRzgDeuM2M
b96sh5KchFfQgJpAFXRBqVmREoy6EJCPaJqvChDGgif9sPqz03QilEaAmtjJIR0GZ3UN5GtukOxZ
ADhslH4vdeqnCG2Z7BZwOokA7M82R25I55tSx23hmm+4bab1Zbg3O7gGW9wX5MES+16rqkSgq8Ig
VLdQFWTCZPViRreJQSu/Vps1xtZYgyn/Pg1PwV4QDpaV0EzKi96MeynIegT2L6NvCZmGbhEH4dqv
wjPSTB/boI89QqmfYqiX/Q/3WpWgzUi5KbE2VWf2gAy6X2QBJBqMyr4JjZspizaPvRIaXhS8COL+
YbNBXaHSiqNblEd2Wkpov/iAefq4kSTNW2YNrsyD9vSHJuMTz3dJd6oVq1ARfCgzHi8oacDnYh4R
wZupXn8ZaH5a1EZNJ/aNBQCZVC/HAblZgTmhYo+3rKMyOZSpvddXD146gcW5hTxXtsSg5n21msmn
YWd6JDzF07kKaPvhbfpbEdVBC2oGNV474T2ry1JJvzMQTyb7Ao1mOynkc5Fdf/nuaVSqmqxhlLPW
/UE3YY3C7+//N+afwNrpbFaR/l/9TMQtYKNcqBEpGvoXQBRA4n4VKv27DX/9MAeFQvt7d2Gp5zHU
vZFH61WTCqxM48s+BE3MROPW2WHBXRsGNYlRh+QKiTwIU04n4ATRGy9KLpvkNFr4a4EBg6qTZeJw
IHy45bNGkS5KM+fPxA2gafodrLK7ZWfPQGxLW1HGsoa51zsUiS7+oivRhjtk4t7FtGwmtQ3s70bL
jZJMFJAj2JoSIUpv5kHJjeXrw/5eyy6N09H00gyz2XGvu0Laa9a9uGLRKTerLHDecX+NMmHGq9KJ
yTNb7QjJDv6KMbDsmYEyRmVLy8j6OZ799WEFSAAA9gFipGPCjCLZoGCyXLJRH/lLSYV+65eBkcZh
WXC7Lu63h/1dR+onavLQ9wgo/K/MKhVBXB++maiuKxiVAxARbxyDhAQhdyPHV/29fnYhwE6syCyH
e0c1xmJnj8CfCRF5d9HkJuCirwDJqUDPZfzWlNa1c9LlhINDG8qXhaEWeQiFrjwm1RwSRuHiOI8p
8JvBxpVg+FmceoizvBQUgw9Roh46YT8S7gt1OE1EP+a9aZsVM4NFJYt82zt/mt59JmO8SqAFPw1Y
hrrbATawr4Tb7xZVNjn+p4Xw6iX8rWj/SG0r8YfUjXCKl1NBuRwiJbeIp2jg1LUp95SXQHlZukTG
0vDhEYJjaB3YYlDSIpRMBZ7ckbVlsmXz1mI/kuqp/PA5TMbmCvW0h9MbsebIQQW0DLUHytPBNGxn
TT2sWGVOZw+1UdQnRYY+YTFCHvKaJrlkw58BKBrAVrESsut4p0kwvKRpQXROS2qRcoSKbYsKwRAh
T3EKS5DraqcFJbjgvk8vU4DJBObAoc08WgtdRZ/JCjPhgTQzTFhBHTJhpY4WeYLxnvDoDcgYA8cs
b9QxZ/U5cv8qxnQ9ZLFl7hZZNxc5m/Eq7PGhDDGo44k76Fs1RopPt8kVJRRNMGgrqAlA6eglwski
c1tT71wD3uHHpeyPzKu/KPvhrvidklAKzjitfLeDdbcaRkexGi/g5WlNjfK09/b59EHKwWl+cV3g
g9Y21xr+8c5g1QCf1ue6fnq/bAOI8LGApxK+00y5NuYmxc7nf2u4G0yngo5egJVJ/HJY1JddVIMw
F8Pjzg5Ci/8108HcNnfr5IP2bShd1qhoYl5nUV54xuCXqH50xXTZwPooN527R4V2URUGyHvvo9R3
FYJEv71mu4Mlw1BNCVNmI34p3Oi3aDq9C3WBtRl3zdnh9grdieg5sATekF7Rm19eOeGdNP3Acf3H
o5Ca+JrSiGALq1ogZhuM5eKnmZnsWUFACXtK9FrbKB5X5oiVvDwKr1CPN3NtU+dYmJ3p5Elcl+Zu
aIetUVR6KmcGSTe0MJ2yRoE0y+bqOo4iItkJ5oGPF6dqRhH6rwb4HfdM/RqwdjpAsFckHYDeCRah
uYwq21UwzV3957F7swWzOb8AlG0PNzhpsz3qbjNOdEQjJPUj8/xWqN0KS6Xm3nuAO1znyo7naslG
JfxmLzW45bzIOlTrPku5IZkrK7AJ7Wvtr19s0cKvpUmufVBqG1uP1MV9JW3Gidc/ez9siy30KQX4
aC3RDx9QpZNeznSGZ5uXeOb7CmWJTWn/NM0N/1m8Nzg1QvO9Ad7LvNYZWpQGQboN25V9XuaTKWtB
MYZqPdjMGA5Mr5acbX82wOurwMOM52//9rAmKC5PyZX/MBS8z3aoVSrEMIwAS7HcBmO9doZzEL2L
3bAf0LG9zmXuyfYFRX1VZYfHouOknSewyv31cSSjSMLcwu5RTz7cIJE9Br6QJujFhv4civGymJEk
Twestc8s4V6ZegorEnTrDsQq+bnRtS+HPvkLM/QidvkpSBVVC0/1qzKWypcpC5CL8q0puQjh92o/
DTY2XNUlFSTrgrdK+6woiKiUs7WD6XOJ0QqaahERvlG7JPIZK2iCmt19sg5HlIRY/03lLGyppjME
FTKhqw8KWBiU6U60R/410umQvuWkZANdB1HT1YMTX2I0fvk+RZpwBfuVJdi7hFJWgWimfVP3miOM
yuz7zj3QndeExLNtMJv05fER25luKFfBFX9LuFBu/GNbCUj5FBPUZQTJBWYEhad+kpGqnaiZXRGf
VNSVkdsuedp3hXkgXOYQJbGELOgt3pbkGyMsnBnHZWNdsbipr5JbrL5XeEfjrlKhTWtR5JAjetOP
EPhLYY1pRg667IH+UfEfARILHaciv/dmcw9GpMlIpYojw1y75KEvPss1ptCgkOE6Ql53U64dQI0Z
N8Li8WgFvjOCUoegRmAhXjRa/6f0VlnAtqWvTLMbZ3t99V95qEiWp44b6h5jVIP2h2rMQufy0KzH
OBORncJsWLIYx1pZTu2rCbOCAejK4+fHEX5uh0uUNLxDM+EInZ3jF7Ouro6AGixUEAqXYu+SWUJB
9I7gvKv9qvmTVnxqK7b1zKqJ4mtdD0xjXO5rqnRc44ljoCSKaQCdKKsaxtoONd3pNb7lpIrUmQ58
FkoyJm4rzAqDb2KyxCLYdLYL/gjD7P5xUwQXs3C5ejuXEqUc1Lz5bBnkxUTvqG12oDQcsS3qT9wk
OliU1sZK9BQOpczyJv73+I/UTsn923MUdHDSfE9GE4kYMY0hVCYtTgV1YwGn1GO8pkXCa65jcFr0
TiEe6IH5jsjD/b11b5y7F8pZIkZKxtSkQ96GQ+OuChlmQBPsY174OxAJIIm2Hw7GKze6UiRdGvQ+
LIXhZ5mZqG13biChke2sg3tSzdI/F2p+jsSsoazK24KrKaagn8bFENDCMTUhzLt9w6Ttwupja6EP
7YpxM2MFuzydq1gJCnKPo9Ny9W3BqHIWmen5G8ygtjqVyRCVlIqFNRVxVEeD3GaR57Kmvy1NotsJ
HypEWP7U2Nl/kkdLLWDT847zbQID6AQIYMEJEKtx1C+ad+tsuTZVF9x9DIXmw9n6LMmy+NdqqizZ
Wcpq4b+h/RGMXCZHeK6LUvEKuQ5sQHLP9SCi0JueO3ED5OXkyeb08lapoz469uhlgW63hk5lY5FM
pJKkq1uGcahV2YeeIvWkuGZGylTpPjP8Fvaj8dJcvbhhcG72ZWA0CsnRLhZNSNnzDAUgL83MU3wU
dn5PtRSrZhSHljcTJj4M9P7l423udL+DaTssbDmhLm2c3PSOUZWe4xFNYznSsCAyWQCLYSsd42cg
9G8kGCNAHZ2ZW2ZEA5L8dXXWn+9adnDV5m8naRA/lBpwPqwQ8BjGOL9B8Qz3z/rJBKlGJuUxrvxl
xIaIZkvHHI1peS+vb4CBmhWw4vAHnOXyhhurhG5m65Vfi2wPNaS69GqA9XJ0F8MTeEUUkgZ9DEYL
Vz4/jqgcCKFqYTRCvsEUHjIDgKv9UzE4WDxA77Dc4NFzGuC4kQrTwmRP7THH+BAE9WCQ0riSXjYQ
bVaGF0412YGk9YcN2DzrvWgU+zZLCLEAWXyyEQFMtuh7nDe9FYC0aSdOgqiclVoWxRRScx8Ykicn
2fAknpXGf/mWNCcGl5wEnsl0WecLZK1GDZvqw0lbY4Cqs7UsBDqe+YHQcVqiKLK4Ar18edy3yH/6
XaqYt6yOiYadMkS2pVwb9rLbYoWe842Adu60ZgWyUbtyi0LY1XfXa+L1UXsBx2NMMWatDOShG681
3vTetEepyxtAiT5XQvDxdZ1sOXuaWLwmmPEtUz4w9W9h6/9mrq8WA+7szPqmyH+t4lbprSorXLGJ
eDOtvGJ44fEXOjz6DD+ZstMlKsdJg4dYVodjg5MAPR4x1jbUbVKnI8ixRPv8pAJiY/3bl6MQexvT
Zax4hkv096n7t+KG88TDtOjzHTXobCxh0iIZTYaQM0vBVbx/tPE7fHQkGKJvZcUTJZ5S3/v2aOjq
Jb3+87ActK79LdSVivoh/tpSb0hk/Is9pWePA0iCnqwlhuUcdjyTmE4AMS8UEmDnutXDaxHNMVsA
7L2qBQaHXVaWZiz5hOc6s5/4ZC1O2ZS8Ucd1wM1SBZPQYBUa7ucby5cPa83SHaWsMrqO4OJFTClE
ZLxGF05k/tJKvOB7E6drFBKU+N/6QhPiGPH8GCsZpTLXxeHtsHgE9ZurMs2hqqTABXPu76AMkiE9
pH2KS8sbiVOlqU0Zs1jtvyPAHPOFYJeBrgYgvk8yO3ecgLpP3EElk4ckvXTk0byBtDbn8A31qVbX
ZQFN311NrDoZ+1S2NtFyMXsRTqt5XW+dLBJjNcWvBGEyWLSeE3VlKvU/MUxp3glNHHbJzvDhDEBZ
A1nw+SP10Y+r8WmhZ2TIzymFegVrPFbRKg642UZnPYq5oCjkWTZmkzf6ZvaRSAubVW70KJCNFRF4
GxjQzulneA1iW9VrW2MrNGyWE036l8zVvFP9i6MjERhjiuOdVELMZcPc4DLCRL1/LTYAItpaFvzK
Xkp5MPKctmGSCqY4YDS8jVb9f3uivsAN3Pr4mNby7TXuX/lp2Jk4y7CJE2ZSG3PuMC0sT2LvNtR4
F01Gpdk0aCDpFHm1gOaTwq2L80bgtKPghacG85AjI6rLkkjEshZGbWAwbEHZiU/VrjJhK/JGu0Gl
x+4Zokf7AszHT7vibpc0hPvDRvGjCFNbLnFrS32H4ApLzC8cIkZ21Cfj8w/LbHWWKFJMzczoJ+ls
YSlEMk9ZDs41h8NoXuQ1tsGjlsV0UxLAYOd2bqxq+hKhHDbudnFJ5V5Xtxn27yx2X2+89o9ksWiv
P43han2AGIdN3KeYlEim1gzwJHLkI3P6+UJqt0oZzg/PyFRVOYz1N99f5y1K2UBcKY4PPuB04B3P
5i5RGPLW3NhFlIn2FbxgUccFzrRKakSkC5zGAg8VhQDW11r2Yv5iv5WkH8E7Ob7eQ59olHIFeRpK
iDKGE3SgdpQgIhk1Gy1+zwqp2HfEKE5NAHEzGB52d+NTCx07xO3D504pIzYpCgQhUro69Z9pwJ81
AJHfG9zyuyYk6hJuZuLanmXWQt9sAqMUEuWoU+Nn9tMgS/mMez7FCmIuSbSHO/JpMlscs7c696Me
o9qsj4u0gnXcWJLK+qAX07sAs/zo0H4jDqyyAPFx5Y8s0L+t1gd/FiINpverq3tl+vZ/7frkdcrY
uyJztYl3S36HhNjfuUt2jDVUyFt1xvBy7AbVvahsg9fOKL1qh3I3ba7ZnvwQiOKoNOYwNkQbiTZy
TDddEwo3RfWzIh93BN0sVP1ARC2WuJSZocbdlkpRTuKz6Py1LICqaMYvBZIsO5+7gnK+ckq+K30J
wtKB6kwd4/vUgn57lr+/lk/JG5qfByL/R7kZIxGGWOeYqC8rGaR0sBk41TG4cQJ2GcGB3kiQsInq
KGDeMvRX1I64TquYVbg+rZxB/yJl0kCIvBvzxW695Y5S2pHipdDS7RjE8SfiV1UAdt+7SdXAFi3V
ojSpsF5DY55PNlVGMOm3aK3YDvlaEZeZgduok3iZRQIPQG2VueNhcSOwCPtIka1ib6c5N/hLOuXT
PlIGpnPCl4KSvE0Z4Ig69Ujug6G0bDlmKoGGlvBGVM9LnefboonXNRn/2QrneWx4lpY0U4sweaCS
aZcC8CuaZbNp8OQksyBEUrqXvIcB1qpVTRvGF1SzQZkeDTKOkrOutOEBMWX8+gw6Nwb5kWge+uXD
nM/XFhXeWv2l8EgII+5doqoNoelPKtb4/rCTteIv+GL4oVkZY03wQWV9jLIY7daPT3onL2neFXTn
QqkQ/L+UzRd8/510cJXsY9VKJJ3gfp/KpXC2dU35Gg4hx1Vo2xhUhPnaVEsM6yYeYSeB4Hw+/VSz
g/bayynrd5IGARddRCVPUHL3jEC5w3b8K7536PdVGYrW7I5+dygVtxemFUH3jYygN9yevK0NXPOt
L+A4gPRrj+YU9raCq7rXONVU/QDEErj8dLIN6M9cM5Z2lk97i/X+utPfbRetJB1tptCMpCYuLN99
F4k7qHAaY8aTDE0ZdSL4FMLXIqenfxgRK05B8pw1CKnk54rIJon7HBpy42iyN6nj7bzGMjiYD9wZ
nByrlmywLeFKVDVkiGV0U4SIu9TF+FQrVYHKyX9Y8o1RkbYSXZjhTj7RNVjyqWAKoNjSVJ1EQGy1
kHzpYgDYgY0tcUUgjDpNDZ5lJSJr3jsBafjU5ps9/RoeefVFP5b9LT6/q+f7UZDEgzLA8RdMtj1U
sjO6XJmCxpbzr9KPTgzqieJJRBxKnY+j1RHXMiaLKEcc21R8mqlBB3+yU5byoZjS3bbUBEIXvVea
UYJDTC3vughZwW47UnVpv035RMBqO36rpBb5LVDmoDSZ+5iOzZgtvrn9No6KYxxPiOzFPx+L3ALI
nS+AFBVwdtqQVQ3hx+OiPmPa1YfVlSfPR8ouPP/W6ISYTELqsaVNTY+qormatrjhQUPt13P6PiiD
y+PUJqbcfPUpqniM3FsTyKs7u3Oz/NXzv8iXRQcrPEDh7J4inh6fskWGsTXNyrcnVK0j9qxN2284
bONWrj5WgzDnfDEqBhICuVGbfVkuFu96y6Ty/wuCG8BH/Gv7YmYuoIgMtaoi1tdQibOOu4oS5hXV
IsedJZdxexVsHTEySCG9sx9Zz6yysFdDDR9oz1YEyR0DFALqtiWZBaxbNZLXkS5tYJvu4F2OVK4A
ywMbyV9bmsjG/j70KX1tAYswgu18TwaDoEtuTotfTv6Ti58ObNuO7LJFBeF57LPAz+P/pMHZ1utn
m9N7+lSceX+dqdc56C5j4VzfMIAYytg6lVsygFiUU/vN01vTNPOQKj9ZqjIMRB0Gr24Z9NyYgQvI
KpfpLqxlmVx03YgKqeQrvhciLqiyIDjkqQpHlQzoFE11ueyn1SSoedPlxibjPdqnfmWRakR7vUgT
zaw07Qaf7gEyfWAlf+oH76HqUl/W5Rf7TaNcSldhIGnCVgm3+xQ4jZ9LZ4lShiptshtqks50i1lD
1JIaxqyZNZDCDLXeDSgZT//vMthgnbWqAtFSWD+Fvq5vOOwzN9v/p6XZ6SjNvJJDMdtV0CWRKqJF
jEBNYOZ6pr/AHgDIm9wBAZbakOhJoOKpR0rIwGkLmmfbmNIbSyqS8zHUilLOEng4193eiieuxlbd
MrB70/VcJnWwwM8z9rFKrl1mwpAkC4bCwYwosJoCPHpFd+82yzZyI9lS8DfPTYSDUEjywYmR0Aos
WRAVHwhLM7lCHErRA3k13RK1r825Gp3I5dqy+W8cBdyKCb53Woz/a3XYJLlUGAprsHdpainPi+zC
6Ei95L0yyJosSTVVUQRUh+SiVY8EdEVp7pzgqvDkPYLx7VcbLOe2gaScwhGXL2K4WsnlgBx7cPnQ
Fqmn3EWa9+k8vzzXcfLFd7nHkwu6VTdtuyVXIcN0MOCHBbXPBu4XppoCj1R4o62CXw699TMG/fdl
O00W584R5fJO4+Yjein/l3dXdphkl8Di3HECcwRfKl9ZZJYXYR5CaMlLRhuP3bytKOak+pQsiTBL
Fc/sFmQbsXAIzk2Kx2erjP9aE+e3RwMlU+h5MbuoZd+/2hLD5yY41SZXG6b+qhtBlxJt/sXy+yn1
hDUdmDskZjTOlrkFXbF6SWZ+Hyw3Z/L7E75vR3IQuJCQAGq2m+MaunR8odq01vCmInN2g+880Ep8
hWM6YXLxdr61Pu8A/26Hv5b/yvw6FyuRAkUw2ypMzzN6L6Z+OPCjQ5Y68gvhkzaZvLjf9C2CK7+5
mEl57nVpmJ18CxsONHHgPTmI8wQwOBT8AyCEkFH9WTri+Sz/+ZCPR9n3suohKeGJu/hK/bR/PL/9
tuD/KkKdx5aru/Ll1b4GbG7k6JrOdB8ClMcgrllQ1CsgSWoO8oefFS4RFQ4s/kYBpwJF9Y0IgSN+
Yx5lRaPBFi0hHG3rEBZMEk5U3vcmZXcg2wjmiy/HSJLNKN6CGTr85wj89DNm6xmQ35CMPWk+SqGA
wTri22FUAbOg3A6rVgXpXELW97Wk3JfNaS/ycU9E3PEETFRreCtc7cdXIgN4BGDkKygM5kXlnyaJ
cUNguckSsSpxtPfsoKoMSDGo3bTGX8yj2tWaL4WGzsvRnph2VxmAWDoc4UVoc8BrcRHoefks/+a6
zzG8mcvrA/J03vDgJ3D+OYDxzag22sl4GNZF1sHBTfbfEzlAvUtt0Q6RzW6dMvvTjiYgCWuXQY/E
4qDVuMuvNTdL6CpMHhHyQ/KO8M5WIP9ywZdpidnQlBSmpOfl/hZvDOf/5egDlGkSBbWnvLnXP49F
ZMIp/diqwAAXxUvko1ih+WbdkvWY4S3gxrVAxNJwk2h0Z/wG7V3OpmDF2hSQct9yEbBF9gmzDtB+
I5FuTqb4R7x2jyNlWfm2BydfAwBCGc3AB8qAiTBI4KZWxtGgsR/u8N9TGR49fxcPnDkHq8Ulmolw
Fpig5OGYomTET3N5ujQBKWN0qz0tZLKJ641ac7Ogn524VDAdnyjCMy4Bdf3pOtmv3EV9pEGrWGBB
+uN5B1sT2nLvKq/flOAKAQt/usghSE+zx2bQ+Rt0JtreyTPl7yI5ByUr1vdq61ep97qRJ6NCm0F2
nNVzCNdCBxJMkYZStKqckCJRl9fiBvvTrP4Xhbfjrlam7DuDQzgCKxxqviNURpAQkfXmcJJ5Ajwz
lMuGInnQN/GvacVK9MsEEUpF9ZUp9b+YEOzClxP3DnJrmP1/vn/Ws/VKvK7EHw30MClVrIm1zf/8
vLaIphLOfI8RZlq4IPFD+toBWPwAHNvjXjZtgN1J1x39UJ+b+2aQmCOAD/aBKBmr1HX0AUY4QpM9
HMkWrPxamlUJWdmMpRoiZVimd2mJBaBcu03BBaMnvemvRSfs05CnimrniL3mHl0DSsPKu83atxQ9
W+9w6zxsHWgoThxlH5QkUU85yKBHBX/t0TR9Agb9ZE3Ht1/Bw4DkmRBZhauwXaixHiliOgsHtTa6
kv1ShGMWGavXdXv6DnMMptTev0x8miHL9Q7mMhvyi+gMpR9EhjdSS2y/s3t4AzmIlkEBVO/0p8l/
LZX3nxnB5CYrMWC13W4Hu6OEn4vKSUBwaI9rw4U/VUwwVMoPLT3b5J1b48meipGpojcroM2xCt8n
DBxzi60tigj5/75rEgotSgFOOGxt9eOpJmnYUjPtCAFXi8NXCiEzbkvHQ+Q3GJAR1/LA4H5Ay9QR
Zl3rU/crHiw/7U2nvTQ6G6z1AqP8W5h3dvqbuwknEJzgRxp3/B1xT9O5sM/D5x1h/tDez9FzEO6L
F3YZO5BKI0SjsI9Aiij8XfHu1mISlkA4nA+QYftQf5WPS9E2tk6hqf6T67D0cTyiBjCWAU9H6ZJw
5686aubSaex+gT5WBfL8MCd0rgkidOHfYQEYZiBTV40mh3YyKAZQWqEuAGqXhcEBhBjsuP3+dpBT
DcXdzZ+uySV4GBcvgN85OfVTT5/Y5wPxKN45r1HyD5HjQyVi6xMvuYEwzTlN2vcyi88CEvv/af7I
ly6ZhLivYpBKGbcmvbijUAwaQkxSsKG86Nwxu2YfTWTw6UR+p2EQfjlRpemzklvW0LqHZEirIggu
kK0vQuHG0At0PuOwileqrEbgU5wso3sz9wwyI0W2SLi2RBmPrw/ptMRCwknlLb9n9v52PrXvYIQ6
18Ee2rw71l73QiauOE5O6TLAkoxaRTQhfMttDqe3mjo+ytdS82o7AbDFlAHbvMBzh/yTSVxsz4Mo
bWVZgsWeVEjzBUOq8t2blg0MCKWBV2+uqdKuNzm6ThOXd0WkNFXNq2LOjKqyv/hiv593HkTqSEnr
6tb+OvbY9v/DxSMe4Qecz/D5I3X8zWw/pLCQuIPUb4/rM7SIwtKlwuQc6ifxa0/OkGn/W4bAYO76
Ou9JI9BrE51yG8GFxHIokKc3vEztsbEDAPQQVo4w6/fMObFuCJsyO42E01y1IX8XIS7yaBBDWxCx
dFoVWS7G5P77NrcUthd0vcsLx+GSg9K7lGgnWxD37a7Dh04lQ8IQt1y2wocp7VnN6CzDPcp/EXFi
QbpQuY4Wpm57XnO1JQ9s/fRKkRG5l44mNSBiR5Ju5RYrth0FPZ7vgdYAsX9mvG+lUugGlaoX6Bim
9gZxMAFQ7htJY7Z92oo5M/G+Qb2FxjcL00Rz8n2hdA5+OooW1lL8Ii+EC8W91RjBd095o60Re8dM
zzo78n3mTnCt6FIedbiC6zpAgEGR1LNBfPnhbBqXnMQd126lxPgmiGtAplgkSSObNW07Sb/7KhfD
EH9kge4Y0VjuTdn2w+nEOxRduzn9TfA8OoUBIr0+0KP/92sO8TpCvq7NKH4Dv1Tb6tT1mGz9eOz6
7bIPioDkInpP0EoXnBaG/MT/gXtfC5NkuFRovtTuU5PB9maYtX+Vxc7FWuv9q7uQJZTQp9ztsbad
t79retUjpWszgYPmDTnyLMovmib2qddyuqDPLrsuX8Ide35Gxbo1050tUJX0QQ00hmczMCVYbUuE
64hfsuLJCXWzIv02cnEFKht2F6vUfWB5QGxMy4D2LUVsvwDzDZnTfPoEW/m3i6elWru11mRPUMhB
nqv4uno/BTZCwqRUo4PYQ53sxo4Bn81sBt4Oido9LW+F/oyPObWX2GLnFRjE9HSv7lG23OYHsjD2
P/dF1+Z/vAZFLAIZUTZl/aB4t8teTVobZ6GWjhzc+MZkLs4HUmMgidRIFD43t2jmAIHpXjFk+5Lg
WI2TVdZ7k+nDCPUM37VXx3G8qnIUYNJIO22JVGkmpICoC43/KBZQ1o88vbM6WUmJtnDsfhMa5ROb
PxfG/C2r7DxFCZbpsO05N1y0xVh21yJfcebJkc8CiuPtKeGpmsM1lwuVlUWRKYOmyMjltfNdCMIQ
kkkVG8XmIc+HUkukeus+1qIXn9UmA0RkM8tcdZDWri8yfjEKJdCzw01V14xVUj9kXHxFuRBdtDRT
waJ88rzulJd4vloxVR5iInnOgUwdYK75broKk4dPH8qeuXhlRS4XuRt5KE4G5JQNWju/nG3QhWqd
onxzKpqjy9WhZ1Hih9FuuuvXBPrK2sj1EVCiiLSEcFX++1kqpDmfqiggMvM5tBASIDEteSvsWNi1
rbxFfu9GG1KuPJzEmC8N0pbBl96zk08RsiUqI4uwjmJnXqlbIzg6di5IushpL+yNdn2euaZYHDlW
8cuytrAOc5HYNsvWQ1XfU7Z1pBQY+evZsnHwqqc9eu3Qx9w7ci1EkVEPtsKBDhCE+Qj0zXe1L94+
j2E0SXNZ9aPKBZp6hCxn8fBDxXCtDr9lU48NcqoQSN8uQ6GkvpZPhgq1opfvCHc4qCf9ds7YvGQm
UqP20MXtuRSQk5/+a2PMa8CfZzecz9Ni94A/bFnSnEMrbRKLe9NOUVQNdAw7j1jT8mUXznvPvTVj
sPRW4W+GneyFcLfcxGlcvt0zdquNgoACxlus5jPQXhzoHgGsUrQLVISx3PZWkkyFkcXw/N5YEusk
yDuccGM0sBHfS58QpuSrztItleKJ09M0xHpXYzzQyPakyRHkSKlooCFLUUp2OmwCvR4pEzEcjyCC
NY93jkfo+y+MGd/bJH2mGtGhEnbIu8jAtsL04q8njRliqMa9EzNSnFiNMdggoQ1dJdVM85ADp47g
Zx6dOuYYR5SQa/RaAiddwtLxoJWRDfShcJBwxjJbhXK3p5WSz/yEiqhKgVTj/M/a5hS27InWa3Rk
B2kGwlEflzKmQd5qGc4Dc+UG/baCa4DAD1l4J/FqupVHSoWqSufI5OTONgeWybdEBJZL4lAxJQnX
oKV6AZv//iUbEKj39L+YKcMU0w/6lA2Sq+LJtDhymX5hN7G+bxGmzApQU1iYk8ud1H7lwxuRa6eE
PfVqtZuQnMMQXEvLUc1Kmh9CROrwpCVv/ZA5UhYyTUUM4Xdb3ALXpY+eQW5R7wuHWzJukoqS4MTA
S40Js7pXCsVwvgCIfi6cBDhbcTBGYZrpfF/5VI4bTc8orsEjP1QlUz+1qGwHS1W+3fM3h1FpIsXh
cr+I+4h+eqfV1+FiGcCNPeTiJjTPZUuwjy30ndp14G9CqODHlyiXn371EoIyuh6L8/2HRz+LAKVy
sE9wDJIYqj1ZVNTB6xuB29A73uCQxYiQQ4/QZY8Tm0XD4aC3Yi6jO3PcQZRS1DJ+flawZlDS3yY9
apMrmoI0qzoFs+CeEVUrkgUWzTARP+Nvo6OL/b9O7TCS0wzJqflL2jWzR/NIpT+p17dVqI1YmiBz
zbTk4PZWq7OP+7dmIcuLEGwtzHgvu/b4AhSeIlKkkJMQ/BRSeDWpRxAGULlStmzaJHdXpUVuyiVP
BC1yBeA3IYCnLQdhi7nzUb/WFuPgkMXdVfByPURFRfHWDV5/q3G4q9UEoT04EWsEXiHXujRdD9Qh
fIlnT+tmaETOeLOGaVuCZZNtPfn1LsWW6ENK11ThOg/iVfCvkQo0J1UwHtay2K1E+qQJAcFGJWgs
/Zv/pvKcrY55pC6SnhYf5FKPIyVsALSxpYm6eG2nfdIZPh2yIrIJz54ypz3x+lOJa/e4vnbGC9GW
Ro0JUKGJjgwIMKEhpUs1JR3of5McuYprB1/4NXF0Mp1yGmtzGuBJdzLH/1uEzwGRC+qvodPDT7Pa
61mfjYHuPmRh96w8dHLnkQeLie/wWWlPN7/WC/WvCq+E5OZ4VtPYxNQxd3nGfybzG/VdXQlmK4Nl
qAKzzZeNCZ0t6CsV3WDmWOV5eGpCAckQQ9awgA08TsD6Dy0UbPsKdYXXvsW1Bk/eeJOgMyBBzakZ
hW6KM7WbuR6DJmYB+zjhRVedVq5lOVF4fJMKVAWhesUccwakXQzg9Ytrf6v9flRmWFsY0zhKJc7C
P/sJE0fs2UXT4ID7Q2f0OsZgBKPKaPyco/n1xfQKLzFOdwqHB1TPSkZ4Mky47OpzCZmTk6MDI92h
KIKW1pMPuMl6ypRZmvzcqXDsP6pwnqvSzbb70xpPphFEt6qnnFSgFj90zISDXeGzvcfDIq2CS/g9
zGCzCzmV9kn7L7zdAMCMLkQOUYt0ItB01C4UT47gYdN2MhoVcGpKOD3YSDdjNYfSVkpu7WmfOerZ
y1zibRgUuhjmApU2uS7ZSkCD86w3Vg4qNfQuEh9brV6D/zKaHval5oyV2mrnzPZE0dV7Nsz13h+2
2Lcj4ROGT5CSpe9yMaC2zHQG6BpVsbyk8+04ApfZl9+gX9v2sk7lI73tJoVDdguYd0VccES6PMWJ
FDAXAUbFWk6ncSrzd6c11Z+v4tWpDKqTjYgL/vVFPMPFwKMJT6U/cct8XhlHz6LMXHz3cQ0Udb3M
8XB8nlWZvQ7/dkO3AUYwpE8jRFN1QDqG5WgcY17/+Djs+Tqvg8IrjIlc5Zo7293+z9cFefDYiXe4
E8J6ctVtiIDto+nuTIj5HwMSsxkDkqIGfImwlmMmkBa0IkqWB6CflAmpCYYI4j+/p5ACw0DhRV6j
laqyUED3TxOUoZ8C/oHjrtT09bUbXNtSKu9JuW5y/lD+VK+zzw153KYGSOUqCkJYq81dHZWWmznL
bASs7UcoyJisYXHDc2Gvq7m43eOUE6NzQ082j7z5rIKA6fsoTvIc4Hb1dQmOJ9PiH/BRfOUZ1Ncu
+mualhbTMGpnnYzNzic+GKu6sok9hZ99SF/4cw+JuS6DMO6nXsKZHFQz096VwNH92oKfwYsts3zR
ehpFcBWP8Gjp6HLAcdDUHOBQPDrCrlSFj16K/eFXqwGuJxycYtGGq5g5ug3Ibmh0wN7+IYq7ARTh
HxEPnSgY8Pz4gwWZyXRbaPtUTUkKc7qr/jlMNyTRZ+5/Np87vxGNmNJKCNRBAD5VtJ9r/LamIjWU
5dIE+0R5+IwO6umB3pxTjwQW/7IiaI1m6/Axg5sFjFExgufSu5YdgJd3kh7s6y4IeN06KdwkuWUa
HF8F4nyQImXg2HWWFrUE7GrXAPGWMZXnHSZeaVRmTPGlff757jNOschlTnn9bi/ZxFxUPMbTgf78
ccBne/RKflsk565/Le3Inv3Sebv1/Xk+m+8Y+ZSMnn4SxjnvbCKVNEINZS8DCG4+IQW5OdvjmqZa
yq9y7avps8pVLMRoMtFODRgaFc2As4YTWiHeOYk+/ouXUh0YbROcoXQGhDUrRSeqG/S49z0xv9Y5
GFLOLbuZOHAWYDQ2gHv6D4R3Lmxkb7AEuK8wOTASXvFPuV8Cnxwxx7/bETJoP5f9nYV3QkuRHS0B
4qREGbZ9z6WX8qaasDkbWHo52u53/oLsYCmOsbF9ALWZEwGtRu+qauOi7LarXksN8O5m2F2jaVj0
86DvgCTBauvBe66wSNWXxeupARYhmcs05Xa+5pMbjxBlk26EIAlCwOdZ+RUVYh+3nzN8ErLVIaRE
odrD1TvP6dcXrK++YwfegqMbThFS72FsAs/YsBHrfe25knpp7TIXrHr8SxlMSeqNQG/2dEQutjsa
2fcPT4pR9DWUD23Tu8ebmGNQpH0558ftaED9gbgL12MM4ADM9t19+tUhTalwWKFqwaMrD4b+XilD
R3M+TqGkfd+wmSyfH58uH4r8WIYwVVyrrd0dR+tiO6ATp7r8RFfaKU5DsSF+uLCPcaPbzaxEWU9z
BY+ofC5FSnjCLdv0PlT4LlbbaqOyteozUQu8eEQROLbszyMD8VeS91ZtFUDRqLcxK2/Sy1pYlAQY
6qP5VntBRSrQrX2GUEnoP7wPPEjD2dFKnpWHUJPrzRpBH5HnGMNPvVRvsSOJjSKfwfT5TVlCQWSn
1yO/9Y9OUZSgdsE68UaUUrs2w6AlwtATvqQ42WmiFXSpG18mcdIZ8imsB8MYZWG4kfgjXZSWfUyX
qKIP9UnGcTM0+0fJTHCxKWN5ZLVqgpPdM+xdFooeeLikvY2ndjLM2TaGxniS2fmw16wHiPC76QNl
AOSz1rWMY5cF2u4ysZ1/otiZTWAoImDfLLzqf6H+50R3UJAx4o328MXaiupWQGTy83OCd9nU+79x
bMkLIdGimu+CYTHUQQzNc4yO7Uc6F5w3eJXoT6OHPGwlhZDJjolUe4aWWnpxRU8IejGkptts5Fxy
hwTX6Wn3oAtnBfYIhgH+nI68f0V4l7KqqqEMebei4ooJU/2g03ynOlLmTCcH9f1ynu1Rcx+lo41F
K/zMkgtG+HZsJefZh1gQ34IXQFujLDxRLXeZBtRmonVp4QnaWdMcUQwNKPJXuWcqIJXzhJ9dtPHV
WFtlXLhnHLlP2C0YNawjk07gWy5gHAuQxb5tfWM3f9oXclv1ZSfTgvGWluCJuEswioq7Ol3gfXzT
y4uWcnXdVZL0S7HCn7sOSbTlZaVJjVLWA73JN+ccftQaeDoJQZ+DPMD7Wd6V3SvDpKSIALId/0hs
Cg+ve/g+mZbmwz/FTfs/mAwvjEt4MAA1hZj6e5jC8y4gwW1u7G+HRtQGfxhX1hFOV0WBLHa85ndv
DLIOIYxkPu+GHUBSrvdppLVrEb5fPPOS1OHkFa1u1Y7CH9zAwrTC7u6zngxBC/zStmMFgqFq3q0i
HK5U8nrtkdpZ4uCUz1Uf1rylTgzUATIWgKR5cJulbaxmc3GE5d/lINbQEZhKV+1hk6qEGlgVQRB/
4RTaZSq3YV4JIZKhzq8Kil51W6Y020JVzqNylIVvUfYO6+mEdMBGOTMcjvKQ33EDWCqt+9SNZaqP
O4rWI2YrNguNnQtaWsQPrUiJ0XCg/Lf7k9SYV7gpX5xua4Utu6ESMlpQYqU2yiQlEcQC3M3ofMoP
4dqN7+7Yt/DTkDX2Szj9IgMdRo/rPLZSZXvi5lmXIqBJvNVEFPFat00+VdSWx3jM1/F1nYA5Eyy0
GH88Hm7AgKQ2a9vD0Ct9PvqUpD8p9JZ0tX6UJme3FPtjtFciNLpNHIETFteBPHoJS0y+XfSJXRrd
I+2HcrlgSeq1W2D8w7fqpG39O8DtWA+olYakoiOxNZc+PfcjyAzVYc7gNNF0CFP5oRf9atTS/PPx
ykLTmN7i5RQ8t+1lOTKXYf4YFXHhkSAjSCvIrdvqGp/kS7oDF5uMDsltTKE2TYpuJS4USed4mzA6
/99kRTgTtf7AIIwADTeOBhC0bftA6VXPOjppQ+jVGS317RMphfq+livtFuslufb1cTLhse/UKEmr
PNbwK+w9qgOvKRlJrtpoJIlNOVViIbc05LIb8B5xEm49phzd9BQPbwIYNnObpENSCUHIwCdBY/l5
LhoT9Gb1iPAEfnc/O6b+3VBbj2XHxZ/0xH5ashtGetwQOa8iBNDj4w2YPNi416kfD7f8o48p9TkK
Yp2NLBh5N5zeqxGiu4yI2C2Ge+xF9OFDLZqkqQGCzAzakO5St+ePbx5coY0ovNnQRW552E2v3WDG
rS9C8YNQlH0a4AYl4JfbJDmExBlNdRrcqCgxGkXtM2O6wqpCM6rCsz+8QKlvsMPXalT8bAG2GX2w
hlI9UJQV3jEWt9AMEuC0//OG5qmWBWS8Ztza8nESpnL9tLq9fQaybpG0ZVOFZGtMzjJ58nfzbU7R
w3GJ0ao/kEVEhTAbD5ggKzF5Y0Q173oIlO4qM81HdAeEgYixjHZ/HonXx90QhTxW8/nkZwDqJ79m
27R1725XVmNeIA8vHM9qciNgTwacmW8IAJwGsl4dM33b42who57mlCVnBDOkOe3mhI1w2+Gl9wP3
Qnj2hYoR9sIu+8shUt72NHMNXuEkMweHp9hUGNGIepkdT+lhz3h2bMLr7rV8GeJyEd1WIZv6q1Ha
06Z54NLXkzJnyJlRs4PSgmUGN9W1t3rm0APSF6aVbfWAWG+6rptPMtUtgNMGSLU0JbCOgJpke35S
lS+OpL6FhwQeaNGmYwnBwGRJHTvj5z1voY9dQ9yVlCXsddhqL6SjvBr4SvYRQWWr5sk65/rjO2ct
dOEoXxMZUNjIg0EC6DXFGgjIUeE7/XqxpwAX1hvbe9QeIKj9iJ0Y4bfXVQgf/azWUF8H5fOVELxX
wtx8GFX39SIskstyWDvDt9FTv44ICSfkuSLHg5EhUp3XdhdoRaVkMILHR3G8mLLwZMABKdn3Igf8
UQ0TQQcs0fV3qP56sqkTIvaTLfC1f3DQvU7I+B8+G2tvegOoCWpb7ic1e/jSHiWJ2i6xwwfeXA5D
dwcL7X6jYmV5jg1Yc7e8hhIOFHKHkq7RtWSbbDrJX+GpKBTAiR8KeHe2I1nnnsUyB+Wh0uK5wWbm
h6CPxI1FDrEMqJCZpFig+pSnjJqS1HDHMn8sR8vrQaqeDPVlx8bekjDALWFHQprYBfxicpyDXJm/
Sqse774g4gqimtXaUChxgPklo0jI7LeErLRzI431/O1eQnAqRXrO3mvCTcIsLkt/icH6YmpndAAQ
tl68PUDunmAy2Id8z2kFrYkyYki2KwpkkrVenGBSoJfHgpy0xKUk8QZRsHjJu8PEXalJks9kgCVd
9uMRWYwXV9GSR7dfCWCNTjIITs1BBnMNMniRY4rs6ZjyfTL5BZfZNNIgFXe1FyPQ9I11LsY5JEja
znK/7h5reFEHIk2qLrAg2Wx64mSNzXdR7f+3SM2df3XyfxNGw9FiAatESwgw3/WvgUH55rTgDZNA
MzXSIDWIqTayk+cxBCgpbexUfp82GDhs6JlBosg0+/6fl4hkGDeholLr2cN+sE9cDZ+amed//MAl
jCas/T0+p41vQsj2ADsrCiuyf5jIpLb2dOcNPqWDOadf1xrn5RD5nR07tWoegYd3EB3p6m5MlE75
0iTByQv1gBbw4K/GUnfiExZ1qHUlC6rBeyI8X0ZAGIel57IX0yWt2dwX76DejOo1eGtmHRR2WafT
PNgzfWdrbyTecXllZ3HYtjfmkyvqvRbYCar9UnDCF1l45QS/m9H30CAhIJYeen4RU1AZRYIcyaDj
ftNZ541rgBL1xVJXMddKYtZLviFTICX+1ROOdNIjvSbhAEokrOeHIe/jNnonHvLBEMPL9IHqbN7e
XNVMLJJxwiO6t0g/uofCFgZRl2dAnycPOAJ6TkrBf3P/nhRCztmD7qN8TiFBzdjYmhz/aP9hoUFT
tbHqq6YAFZgx6RxGpZgTRW9GvmUBHbBKGshUZgD+6Zod9wpcwAKVR4WgGjaYwHiv3hyNJCsycKqD
uyvOjXVdM6W9z9opZiOe9KrwUaLukEr2koLdAktby+OvaYXNehwZKBXLIBF4fB4s5Tbhs+u5ifTS
4Tbe0yxJbfUkbg2SiSQ9wNaxCpReafBxVmUYikijwrR0eStf9icbHKS5MgqZIcJoTvU1JQSJUw1P
2UqO1YorWVQIgi6qhYZo9Bl67hGslLRAgzM8SedEK4dy/2XEa64oQjHx3n8cCTArQgcMc5NzeTXG
VVRa5KKGdbpLvySVtuQO9ucCg8zt+xMhAvI84a69buzEQwufnF8RsN3pVngOYJwld/U/HY2JOehu
m720ht55JpNOHRskcYnJqaPwz8ofWPg+M8nTPAkl9l8k9wzOWmitBqvoTU/t2qFUqT9ShmZE5890
lD3LAeqAiiKcg8sFj91nZrHQuOmUkP8qlEYJFhcL8n03N7zWH54xoOnKkSSW4SeW0lf/LQoW1yPL
Xl+HW+DUszK4caaeQS2bs5vqF0YuIUB7ORhJfdsQjuAEVbThqU2kkNOiWcu2jyEbQV1edUml4U9R
d616JY1PvFgJEGhPzklQiGk6qKd6BXLexmFTwnq/CGEul0QTuUDiVRT4yT/BZhwdqEq9EZKzuVGz
PMCUU/JzBdrMKEyQBiSpyOrDKTCeutm0ADSWUfoxxC2SmvKU0+qEMK7zWpfFr4+e1k6wUzhiwbmg
I2V1Dz7zAbeW+8ty5Fz7y3sXbD+4xY6MfYY7eMFEDI9b0pOgTTtPwdPDq1uQsafSwOMsp4udbbf+
zrF+R9gBqr5z2Ls5bDOSg9G6nNmOYFWw8K1zIQ/OpIBaUaHp/xGdkLslzNEaEFM7F3PelaxTiwEK
8KMULlw6h31UyAT1B9YeRMDSt/2Rlk9L/4awgbsyBgUhpAXKQgFLaqb0RgOAOj/qyUcMCIc0gvy+
75KPEWB5X4YgdQttgDOLsk4Hw2L2LoKwqOlLObg7v7agGZ9qQvfLls2bbpEiMsH6TJXPcTbgrCxY
ZysU8ozuRVYuwRf1W+pXCQ97As1qTcI6mL8MLE+BT6E7ucjegTJaVWQ409jxT0VyEAeNob5vaBqM
zpULmtdqgj4Sdrmh6uHc7dezs8EUM/uPMEByLxWBKUgIdsYNWwJXeNVuemYeczLKnBcIxkc54u94
87vGE7rBZZ7hKXDgdqr5fpDjO4ThYd2B4aVXsLypz8RDC7Pz3terO/Lud4sfbNrI9uP2GU3oYDfE
qwyX0o5C+TPo3hi1TK0nRT7WRdMl+xhmF5KU/0Ff0NEWWkNpTx8F7eRxDxAskcWlIMMbu9nDJQtB
4NpOBIj6AwvUYkq+TxWCQu4W7a+CU2ibXhg9N7i9qMfpwRFr/15WMq9ka1lZdasBMRvCRR92ZH+a
8O4ak9kN+ultU8HC/0CTavsguLjOi5s6nC1Op1dd18DomZwjdKyl5PezSQ+6mSUP6pIL4ilr19F8
AlVB7V/V/fpDFkvDZBaaR10etlgCH2baNUKybmqpOkEQCKbn7BNDQFInAGaAV+PDfxJSPcA+gXyz
MKsDapGdJgJEwBc/+FrS8rc0YOXEYmFag+aRMODQi0MIui85o47Mtn/+U8aoQVw3azNA0JhZACQR
KtFcQSbQzogjWv4h6fE7bIIYtxkmjYDOqkglT3VW4lF7CMh1ZyFfwIZmy84x6defisJTIi7+FhkI
fs3FVgC7j/ssyjAA+mMAZ6JfA7t3A5WfKbps3cMc/erWAoynjJgY+eUFEUmF2P69NQ+3nnduIS+K
hnbznUEba1SigfP1tWR4EapSLAbrXlrsbs4WVy+MgcpqqyqMdP1QifhQqnZNo7dEZ/cbmGwK2G5+
JV07qScqzNggGq1VEVjdYJwOE4jS//rmdKq8pJvQgbcl7rE0KIT15rYPF1xbG/2V8ZosbAh1nghd
NYJ7XcCZlCGyW1pULU5Rtn7UIweTOh21Nw2Pk1a1v8PM+ued1Xs3Wo5lYw65SIdCah/TWA1QCy+p
a9EkUnVMTIUIowgaJOGFqiFyCdItQmkOpo1nO+uOcD9Mmo7vgvSqrQt4mPat2NCjN3XzuFs9hHZl
tyP+wn+2AK2cP8Z18D5hVesD7Lu6mZruyozTRGe0CngPZ1CMihb0B6ijXsxsE9UQnbqgPrTLS1+S
j6UMFqWn/jnt75p2dFPAnBYAO38etxdyMCGadWVgZBXQZ3ClamVtqs7eXyqHL2nBVfmbWfUQmP/r
if4ASLVB9+LAABAQDGiieSdh9N4mDlyF7aZpBFP0jtWWm/U2L2vTWXtFnF06stY59Bp0aB8xyjEs
7jQ1cXG9AccqZShXYbbBMXJtcuOMFNVckO4pyR5vV15YeBkdZso0Z2eqn2w7KO8+N+10DHE8+JMj
LuuBfczIGYwjNqXdIaj6DRIpMxXKwv7WhAUxoaiXwQ7J4Q4MB0BKkyqXGtCBf/mIC9B872r0ebY5
qYronlNY5LPic2Ghwyv39H6wnWg+jzwBhEtN14L7XGy4a+GdhKlM18ua6hyud3TUrlyRYDuJrgec
NjNt8c0HUueGWcZ+HBHrCsQxi1GyN1TrePMlLxiXf8x2HaaPTKofntHWBSvRMVjYDODs+c44xoRC
SwAH5alc01eMPoSSIC2cjMmYuqu9qAD73kPGC5TXAmW27vjjcsTgZ54JMTYztgYMM7LWrsLdQ9Jx
n3QCPIedDWzffSjZeceRGkscpf6/sZh2QFELqrlPt0lrROj8bUsTtucNEZSHbJfuN0lPiDhFTf1k
HOTDUSR5vo+icT65QQ0uLSP3QIRYXv3H2FLLZelHbSfjFaLyUKsPPLKjhzCgFF0P7SYXpjfiLngz
0yqHCGSIXHVL2oybmHbVXlBS9MMdK+5WLvgaf9SrcnB/du3qCcp18rjAYtYGmNIJCZITnIGvQdDl
bRMRZk3CnW2jE1PZbSuVmzosCi93d0gERYoKNh22grClZuaudfJ86kKCZ3yXbIJ2+hWmq/tMYZLt
xsx6vA0p2QZLa8VSlepLoUeTAw+IoNxgflO3Wu8R0m4sicnZqaQgCQQRPsW8tUmt3tfCsth3jJDI
oFIwQTsIJMA+anCPsdh0uG00QHT/QM0z2myM1bBCX/8d0blao3SD7/v2p/xBeaTOtwqeMejATIq5
JvruNKXg0qrH2CHKsjXu+883M6da05b15sgYcV4PYbyJAO0BBavZG8z2m77Nr4l7BLWGvvFrvQDZ
PEBp9nl7JTGFuYK2Nx6crOTebuLR0ROqL3O4Sa4G2FfkKc+d0qDmFEZPRlOPRLLsGpFAuAR09D6F
yZ3YfnTuZYtLRiyPMRKU7HLyGjs+8+PhsIaCiQxjVEt0oas29imjy3SLtmEOMaipQJbhwJ8gom7z
69R9Knd9PoCYORfA0+UxSo/KHs6X2Edhk6Op9vPa8NrNiy6mdMfBq7Yy4PkzR3pJgQINrU0Ytcma
u8s+PFmfWE0T12wWSq8Ay1RkJnrte9PbQGRHWZQYhNRoZfRbVJ7ySeI8yy3vqOSvS6+6ceaB6vrR
7CTetmAoD+PHuOivbOuOZK+oMmpCPbAvu28ElWgBwoMSbWXHkLJ5B+FyKyuftbPQbPRp8IQZDZ3C
lTy4r7RW+BqnRRljmE06j4XmmRg7GSIDaRU4dUMOkfCJpny+fHf2BwFOMxz3fdhX1ycP9qUvSwh9
iS98+X6mbuvvGjLHWERPatUsBO12O7b0PtFlPKNZcbPHpdUbCFOAB/SUWPq8bJ3TmqoS+jpFoAAe
n316IpgbjOLYjpnVDBD1Eq2aEW+ojGuUrwFanDjCAZi73tjqWhoSVv8A3o/LGOZO2yvwoXibhCOU
PlMRfa0sRQToWtHB7g3d3Kb3o2R0vr7++HXs/nvbNlwjX0CWregWK+aNRE142kRj7iOfHmPIhltJ
vXf9p2dgemzUSevS8kI6sNn16/v2ZMC8E4POe11WgULtTy7j92yIkeiWUbqhdd/nJcIWZIDUlrfK
6g4jNupguFM7hbEhvUvyumbbfJ0lzRzIOVmLW9Hasu+WWa/oJn3/2HImMTmFJs9gapVWYBAZu073
aehNnaj1QLAIsPJP8Fo1B2cJkFOVI9dpLGH2JCRpRMHRMvvpwWM/JslEqyCK1ZlHYw0YWMRs2onc
Wc4ejrtuZGrVEsDiBZbZjeoD5EvFwnIbloYqz5MrZ8kI1OYKPD/PdUdrqpzhCjjeN9krCjRGUn86
GjRrKk53BAntk03SQorySIGYlUGdHssoiySXfW99AX3ik1KVSHLR9dchTT7CtQ4DC3scHcBfl6Eb
XEIPO17PaRjzdkIjjKX79UlKjKchASAMJ3dsobRbFXivlwStDtv5Df2uKauVbO+GCyZ3Hkuup4Y7
BFUIgRBhAz75+Oe3RaAN2uMR2oDy/e509rQuDWv3ImsmvKI8Fx/CmGyqrT20jyBdFWixgizYwlCr
q6OQaqjXLPVruuBqEZtQ85NNsQZulp+FmGpsbUgpPsqurYRfT2Qmel/BpviH8Y3Lc+RbISCrpzYa
uFRcLl1yovfoqlCz43LWXwGQSJcMN3ojU7kZ0XdZ6Wg2LO9iyXvAjS5oF6Ai3ofcS5hzeoNp05NA
1LF/yyAMDIcobllMuyyVmN+33bFdIFvP7XlmcU0hBXWbsPTN/oDcvBSlAThVHTuyXB/8gowmHC98
/NLN4Bdr2lMkiVvi9JNLIW4/KEl2FXS7I3EVXchBslgDKiDSip9IWA7/WqIBmJ/vzLVzeBiKb2WK
F4Imm5rmOzle4jjDwWrbePQ60F+Y6RFxff3fEzLILPg5HBrDZTY8I7rFTq0yfh/uz8D7uVbJ8YTQ
Q5reDf8K374qlFMQ5zJM+Paxy8Sd32SsNhwMmdqD1Eb+1bUnlcLeScmM/KwF/jE+a6+K2o+vt69T
hXIUtCuP5TlMMbQVyNdFySFCnoOnAOV3FL6HpW+f7yt2dX/RyrYZrHUGMcVL5kQkQctTv1dV6vCk
Bo4rF79LBfnCY0nDugtkrBgMggkQ4jbyp62W8ZvukDGdJdQhEXJ31nAwMg9teitmj3DXxOWeBj3y
r8B2P674G4NU1mkb740Hiq96L73nKybJPFuLYY506+QdF3JkcP4bba1yMNmdI2p8au5AJOh21fE1
/9t7Ir5iT7anY0Yd21GxRE+EEev0GtmFSf8j4oHLfgwmgyZHLhDaGdOylvmSoCbkYeKyYDi7rxKL
uOVePuXGCXhb+UbT6qjKEUXQ4396MlhlKGBnc1Nt5pgLF9LrYEzuLgCVdkuq5G8d4Prn3azbkaQq
hh0yIElYkYGPddi7YYVdnPluY8y2mB2k+DYA95HdvpttL3bmzITq0DNNgfvOEjbSVnqfk1Y1BUKh
DZdY8BtDaIZhgn1bwSN/kU7mkwBUBPBqmhHFc8bNOFYsc6TUIRCZn/RsUEA+HsInJVC2ciGXvLsB
T8nV/VRq5mV2Es8WV6TjknpwP/yrmK66refY6k3Agq6pDdyaJTp/33q1vWV0lgg3h4FvNcm0GKrV
nBGJnxbD4DZBuF8HdT90+Fp5U1F1tCAiLkOeaj7HgXx3mAZ0s5Brw5BZE0Ux81mO3aKtiZsPK8dm
EYnsEzm8lL2suQoSLbh7dSBDSgOqIySRaMdqfu2ESjptrvZhlOvy5hjXduiWiNXa5kljp6ly0WQ4
cYRpsBnI4LosrXGqqbJqZiP9fusYAPjP/y+jsZovgYxHxYr0JoqBkdKMQPwN6SgPnKpp4ld/R9oC
rVYlYUGxaz+ENDhZ6oUVu4qaj83JV6puArGvaVPT6JX6sG6xk2sjhN72Iz75/QzS+QoW5ZI1evO3
lpuNnWaGKIUsxEAbv73u9IQGspUGaFnDVImxjl6sTCsDFUyagGcK3z7S/YkgHldmokCmJnU5TyV6
Z4kRXOlZxs6jwhjjBcdVGyFXvph//93xudYxOMmVPUTz9nwqCOr1OjLM9kKZEQx7fNlwwPUUV2FJ
ttlYTIxFilRNjDA1xh9XoFCZ9WN9rf2WJ6ZJ7mzrMt0nGOgzwx+bKCKtyZeHeQD5nRjYKLW/QjUS
3Bqw7N8Wtynvv3y2Xo/PpyMoexJNF7+SuGfbvjdyY6fxjIjP84QQkgH382G51WfpmePc6681ZF0J
VDf5uIxQQsRP6PG2A+X1DV0zozAbVuYtjCnd06WiD0KDxtF0uchIPdfSn5FxnwjBaIt4uvtWGbSl
PT30ZZzfdUEGnyLJE0imlJXUwKZ/DJmxqXIXURKjF8GU7fgt3uP0nyWdTZHpSTAPbv8evQ1z2qxx
XwvhzxaUk1hn9agZe5W+kwWrRCJ14Jmfx6GXPwZyUjzroWRXN73kyt2jp+VA5y1CKjAllMF0JEXr
JkR/t00rA+j+gIPVicUfxXIG/qG8qxWwQYDLZSsDEu/Cpz2rWjN8xsX3XItUq6hZUBHApdVhel9R
XdchcoGvPD1DeJMKIWJrI7KW5PEO9UBr+elue90CWvtd/aJ3BIjBDO9zvRidLX26wHd7xnd8b3pF
tAcEOip9nwoX/v0czEVCr1O96G2OB15v7PhqTmNmAXhLX5pwOBKrpC3qSlvw1VTLpEb4M+Yf/FKg
GRabUcvN9ptuWM1rrB7JZjuJ1I5VZsxh5EdpYKWNobO3OqkG6f0bm2O8aVLuA12sbCSS/Khfsa1K
mdHH8Ag4anFVUPVid3/QwriIYEEqzIl+rPeZy3eNKv1EweQEygbk5U/tjVGPw65h+9KaVoLm+kj+
9oAPnAxDZ2I2LDnonP9u0nbrQlQLIr0oGZ7n7C8QtG23CkMpJWmFJz8qAbhImJ6BL7DB6Btjg3eP
4dnfaBadn/E+TA+Jhv3XkXzJDhGmi6bNm2zRknWQMqG8EyN1IHX4wJLXSDK1yRNIsBKqSTbWT7ln
esqU1MVOER5PiKUqjusDYLHl1Q+pz4fBVsJRGXr6p9UMKEr2YQMsVNHIodZGmYKPezaQX/+GANnA
ZyMC4LxfiCySQbbrw3CqH6Ca62IZ35bjfRI/n6gQFScjA2cFUqOPsHEwN/VMIE6Wxhw69qWJvI7K
U5AfJN7uy2JNaorqAtNBaQi18/QzLeHriQqEbjkL0cD3EHFz+hLkUyQcHEjGTuy/xoXYriMWvyLY
+ANUALzkRt5YUfwZGsu0/ZrVf3fC9JiP5+r2rTIYTRvJ1Wa+K6n3dAI3T8zxV9Rap9WeNuToOhMA
Q6r+OeIeU6qjaukmd864VuCFB0dvie4MY1YfsIo7u7SBoN+uP6zZyVFowpZy81dVtz38tv91Tbpg
FQAhMn+RHeWxkxn3sX+5K2ImM0ifg4HaUOHbNDIHGZ0KG6aLSxA5xmyciHTWyeKIkI0x6SLVNj5B
2SSit3Z3bhMmPNPVVkJ0syKoa6NONBxLYWO5rLfsPb9IC5Erei9KK83EofI+99Ac41EB4MvXUVaU
+0/WScaiwH0cMfsM/Epyb+BCtGFtTjzD7oTBACMMOuCKJXcqpu0s9W+ck3PcA3PPNCpEYOrJB52/
6z5vdtdQWTnoJcROEku2VLTn/9jAvP6Xpf91Iqf2N3AA0PDlKaJ7UNs/IjMm6Ds5gPaYA34Rf7nt
4cQJ0sktMIT7buUPUpU/CMhgjsQB6ko/LlNbCiLAAwa5xd/pLemrSp8OD0Zt7VJKQNFSFQHwJLkj
27Nyh6TTaApN1P27VbkAsI8/Yl4VHSRf9ubsMnsjVTF4OSZxcNDhNdA5aDSdwrD2cs9qYbJG4hKw
Zf1r+GXa1oPq3YX6Sbn6W9GtB/7n6PXJm9INl/faoQawsHSvZhqcbXfge+CSXPeWcEC6IZvly9XB
+J39+OxwSwIMkL9Iw5zLD+EqinGfUCkGgXfW0JtXBuHbDdsCWTonnAaFbmD1MyVpBxqN0fx+JwJB
ORIjaL13upJNNr4XlOq1eXVyQOZlUBGOLtffrDVUPTXB6E3I+z7PZpAL/F7JblZW+hYMM74ovOul
1OmZIZ2XfRHyOwFMKI9OW9EA/Rqc8PZY9IBNnDOOZigbX5ULWYNvAWfX3VMQj8rL82kNJ5yT9IAE
VxQ2aTyFzU4qKGxFdVWPKSAP46o9fZ/cc+Ql1gznhGuOIEn1QrlyTcEnoWzwJQHIosg5gEyZ5HtX
gMAgIuKwl42X8WTMB9vPTfBcLjl5wNWLrjdlhyyt4ynENWz6cLfgvftrXHiCoKx0bXpULCjwr+G5
i30yqmVRKE221wppqb473tVKAFAzlx7Dr4WgrcOExcB+orhuMvPXx8uPZjnQGl+akNxpYU5q89fp
MNPnfhZrIRuw4LKRBXnczaKzn08LzWe3FgmyTVqT0Jwtcfa6yb3rIWQgw2LloC+1YVvouxIWH/0A
Ca26lDJPSmRWBASTuUgqHNQxjURDyCh1yMn7xqY7XxaJfP3Nz29GqqOp4erjM+pGICpgZj3XLoGW
YAv6yIzFwnF1uZg64y5KseN7xYCAqF90y876f+vOQoqOQHosd9Kn/cJHluz4bsyOn9Vp1BX+rL4r
vcxkVZ4wEyy6lvmEu1FrN0+Ilx/uGcsppUU0Orni3S27RkJETEv9TwUAyr5xp3tkutdfNtM0QFED
ouebzCnQqCh7pZVlf+oicv4qOBPMSJK0tNnJvfnlV+Jg++tRch3ZIauaf3mwPk3igBEdTf2RyCsS
RWHpQtfV5NzhBFrohpfKrSCpJ2fNSh77wsp+HYHINVZcAatFnstXscxyKqvQ87+gBiFdRzp7dmqX
l1Qv1mHGM8PbIA3mfTnvWJmxq71vuur73tx70Tn5iTv/yshBJ4oh+FQ+ISfVSrKbUewQ0319DaP1
RZSUJ/UhxLpUC6bcaQxaQd7eg3g5mAYUo3s4SmnjQRi/cCumStYZMUAP70Zivbqk9+fnZajcJ78Y
oXwITRCvdPdO8MFQGaoMyLJtpReMMaDU7iJpXL92hE7PjaHgbwtYpGyDnk+EQc/V0deGiK3l8yRl
OJ+P0qhdmcurbX4a0b8kxwGEY5q9sBEZUCsSeOUW3hTFm5Lm0AR2igfv3Ow1HseKIQD5frVsWAGC
jqNJIdTHWXTlpyNbVLtTBABPQSNYJh02Fl+IWM3pgsfOibmBZLvRbnJEtM+iCnGxuf71IeuqqZX7
Jjb7wyWY8nfjV1Mt5q0ATv7hfqEVACk8tI+ET1MIoTLvxvPOkzBGSfAzT9fxqTn/tNGPg6c2Gtcn
Y6rS6vYNjOaAIIRgYzsSh3+qeqO+UJocnfd8IeWEs5DmyPdbAa5VGlrOC8ZEBundyd2PyjlfJnJR
cAuUlV7amaVY2BgCdraadW530PYEIT3gcoVSDgLo09q47Xi0va8xbipTEZv0hJEz8fIDfD9utfRW
+QhHWKj2UdjRXsR28AdMxoslBzNPvBNcjZsW/XkHVMp+tfFGdfCIM4Aaq5w/vKkdH3ia2U1SHTD2
AnFdX2MNp6OFJauiIwYZJGI7sHegxzzhH29LY14nBWNuetQHY71tjxig9NzrkJ4KQzXCVy03IvWS
YCJFbrSb2DoQKHR56ZGsSmTzPVqoIJ2KsrXtpRpqV1M8lilXU0F/b+9Gd6qfDM0cgn75MOXxN5iw
Bp8h8YDIzmcxV64iNB7M47Rs+YG6OzO/z0RcLeFyDiDpyW0gM8qsWhyepg0YUEDlrX9QwV4cgofu
C3G4D1wqn6toSyhAFmKfZZMTdH3Fmj6eV91VVnN2lPiPNPnRR4V29G5Ko7cG+aXuC3nSYrKswVBY
k7tHCYsNXFlN06gxwUdl4Ez9Dh/zakIRCuyWf8+juaQWPzt1hwACg0MKq/drP4A/gOnne1N9rJv1
pWEwST6VLRHJYxjN/l9L2xSQ3ISJx+5G0rWXLM3z9nYFfqxdLzV/WEDX4iM6LB3n4hcBboi7nDzW
FYavGZy7xItq1I5HWGSPQxL2krVqpz9VVSaNPiiUMvsd46s/A0HQfeT8muW6Nfl4+OwiBjMsbg6f
baiuS1e4OVKIUXu5P69gj1o/35iZycdBEtb6Y5MA5SI2wyjrJ2V1xcMz/a+34IAoQO5SP+ddpY8w
m4MIV8gmab7l+ZR/8X7Aj/7U5NNHLVOJFmoEO/z8JgOdJ8N+GdrfZ1mereD60DUHRFikZGM4Irum
oX2Pq2yOrdtFCY4x7bGh8u3bgag7VhkSSffcCj/3GQJN39msEQiwHT6m6nPJ9Y6hObLzsYjw0hRD
d0fdEfn9ojSQftkWWN+GVyQQ/WfFsp4kRl3+pu+Grjb7N/16rC9rdIVDwvrMS6Zd0i8w+r9Nbolv
OZJzNEBrCHU/rxNkvy6O1w3AqhmmjcltfJ4VjWiHyEsniGxBeofwVXLoboU7jH03hIi9sEasB/Ms
UTy3BHvhI70+ACgfXi40b7vpt4yEwmxnuq2ji0Q1ylH5y1zX7PGHE8RLVgsHmr0HJS59YFWZRzx1
+dE8suc9rQhX9pKA5aqoIDsxdkqMh2WBws4aeiA4kdon/Q5Wa1GE7BxNHICgCtf276cBqFkGxisn
ptqb0AORvby7F0KNvWAbTd854ZodiEwz59tE6MbIrnwQPi0w172bsOhf6bFKXdVZ3mq2ypgbLU7N
/cbTPJL2//oyCD1wHgWEWstn3TVfUT4J+dTcK+xjHpXYZ0bPrxmAP8ioQVsdjvgb3pQsoFH74quk
m9FoUsEPxKEDyFtvfhppyy85LKj4zLcOM1eOodqsLFgwe9Xqjf/nQb12RTVUPJkd1r1h0kmnsEUW
jcpQuZcTrsDKHMG9K52v7A5J9X4f9GLx3v5XrhqxwRdLkiToH6Jh1JDi1a/pdsMpop4Zd75KOq7F
Y5U8dVHP26pNdIpmdI3h/kZTA3FLeTzplaXa2Rh+LRxMnZvhvnv4drF1780o08oAmcBXUCbu6rFt
ObpdAXoRpi77ZhtblmBw5ia/Yz3qKjbh9TpBu+85ilnNQQkPA82BhZo7L51C8SPJAMT4Nxvq1i33
nv/8DJef6yvCOtixjF7M8qhJI3OprC9j10GTZYWM7ZgugImhrpXfUd+y/xGE0dhLgiHMt9bEDJ/s
znQLTDpqK6Y22QVeOSm4z+WPydMg60+jtiq0HPDqMeh8NnOr4xJT/7TURhh78gdMSFpHrocnAMhB
kOeRjKFN69WxZEZ/5E75EmgtOucLHTF7Dc0o6s+pCo8ZKNAGWuCU0QnbgTI7U7vs6IjP63jii5ap
O8MQkGSke2iLjX4qJMZED6Uws0uyTOn1Mf+l59OnlfAYHRpD0rd13qHr6XXwSPqccyBh5cJf/5+L
Fh5mMZ4nk8pjA01yNnVRG7JZqv9LrJJ3BU0GHHHpj6ruoVul9cMffB9uNv4yXqNzvdOM0MmAN1Xi
YfA3B6vAYX36sHMX/Q0mBK4D1W8S/RHC4eI1tLop3HO6Lgw/BPDjsyMGlZguk3PdRv4jQVPW6DpE
CQxtn5O693q6Gi1D6Xay25XuP6RyHd6AbLkI2eDTjamAhVd9F5rjOLpDMwv2pZ2tnNgn+n1m/0r1
N6wCD0F5mGduSYUMFLdHOO4mHLfCU7UWSbEMbaH7R/MYq8nawcVYEmr/GpwgKCK7IcfTicdRL6bN
iPPDZUVAu/6tVpQ6Gr2u6iPqCOOSrIWyiBv9NZIGbgDJfXlpLvd0NGLc3SLZ4DpiMXh3zqkj+d8Z
v9SAYIgz3KisFZUM1U0mEdscog1FHe0e8T+TgPEaaTeWzkQShdG8a4tlmw3KX60e4cSMSZIEEkmK
tiUsDdMhP2xNsIhwLZ0bKdih/FnOEAWJ7BlAb3S7PdcuUdCEKW+IdFbFBBMJu3IzxRfWbbfZzP4L
588hTHdMJZeCWsIaK+gypPG499GSg1VTqmHJG4pwC+nwF4QB5WOYOx00Pdy4TlCuFnfUgY54GnqT
k8kndWtR7XEUEfKjpSHVzYOJBAN79CTkZKgRVkHmxXFtrh8oP9hjTI4sbD1IwgiwaJ72ANnrIGbH
gRYzfzu/LtAkiGq0sK0wG4vv0c791N8ncI7NGJLPq6dT/bq+CLucCxPjK7U0UDiykG6AxYHr1oZh
ObyzxZ3oeuP0JwMowD7paDsL2brSerF/pV+oCxjB/rbi0wnjKm0D/tneILlofMUsCYdZCv/Ch/c2
pURMWhKtx47Ld5/Hvm92SOpvpJ2oh5+Tiruj2h8B5qmHzJUPf0iZYgA4iXIwmZiBMeNajbCCX+GA
JO/GhVXqPro9fmoxrX/GdoRll4BSOIbYOdAk1TYzGwAZx9gSaE/qrLLxl3cFtgmYFtg9TH1Y5dEz
TVtT5VEQ0iBRRA2dEc7hLSCUxAAcOpV/kdfeGsmaSBvDw5OcCODO9zlt8XI4BJUxt4sNssuwp+pa
Fced9KFOfSVOQ/JLCgyiJcT8v5iPdBA1VqcqKdKB1W7J1xlg8rxepcsvfTWbHY3iTFhqbTy4jHwS
O5sVoXFRP1airiwMyhod13I/NCx5a+gTnS734heYztB3luj2LVknlIY7MkpEJuFk8SZkRpdooRPU
xkPhSlFuVAOdEP4w94GKqE2sX+/BTnMm9X/a0p5bUI+PnDx+nw+ZlsQDTuZ7/dPQln3imHiTZgCm
A2gxi6NyLI3OTq+US50eVjeiuv1gh5HmIJ1s4pC7yLj4+7FasW+OouC9eTqPYaCZS2LPI1ic22ic
Yc+NchZ4TvF/h01ROv0KiK0COlEJ1KzAis2FqvDcN4Em760xIudg5FGGxpcE5DZGVZ1TUKJbuS4q
GsM0SMDhdGBoPBJ2aac3g2TBrCHZP9O+Pp5SSQLqez1MGawwVCOaMMZbJ9ylDhtR1rjdhnW4eO3D
g+ZurtyxYZ8YvkEdohUbXWs2+NfzkSU2hhhV9MWKZr/iScSpjkMf4ZSofFeVT7t/akekrN/TLebs
a4KPaMu6WXvMvpo3Ft6kEwynqFr9sVm0YDd31Upx8LYCK23ZxW3m+ijFH4LArOBgvXU4mQscooV6
L0wUmBRORmcfCTmd/Hhpo6gsIzms6uKhdY0qMbwDF1dgVfiPgkgWZEo6A0XVIQNCQ0boRYCiLLQi
JobPcIeCFxIz6Re92kcek70IMtES9Uz/BWooiOuem+gpCxL/iyRsCNdeSTYkZHvzxJauJS+NHuCt
8Lh/XbbZ1aDCa085oJtPxDsdkuJWSBP60u1jxYs2KJIfcqSdH5xUPdOIssuASXt941yvKHNdG6ZM
HaMBAvSuc7Rvuwy01ZVtGNsDg33fIOrsa1qqIB7Fk5c6SIXrGSlwGy/FE8pCf3k4SBH8cbY6NK1k
QZNYxA3YErNefGL4JSRMno1GnStWePS20eZtI+DnRD55Od/VkfSDP9NSenEf6BDn/VfOM0qW+9Gl
ctltH3wIAwLgVbrKKFQb5gOlNGxwVUK7WoXGyGM1JxQDhL8MrdeMhVOFcnEz01f5holpE4OVI1Ly
M8LqJBJP9/YUdenq0ykz9GSnM2mlWrOJSn1x+wu2GFvE/v4GuvWVihs6PJmD30GLuGZBrnbPec1i
WkpyImRyRNfaTKyGx6BlLm/+6IMNSwWYD2auNo1AJhz5XmO964Dk2pm9plXQPLzCHDsCeE3am8wz
/kTSAiCNYp8OfPWy3xTnoESrAq+jghwomHE0WKS5vMNZfKxW/3LNOPQxeHKRoX9Zo2w1WCZvtjgL
IlubSGmi54I+VG4YMVTuCUvoc9rfGqvv/v1mu1ys3ZAH3GCSrGm/v4Qf0iBka6R5mpKlEjdtbw4S
rqxiISXm2mWgbA0nH1Hofnkm/wB3sKrqQjrp/VDXfvyfYmhMG9OF0umB9zG9WO6yZCFvp1QyB3mO
87zp/yZC4VrglAHNsFH4heT11uapFv2W1qlM8vSK9A82NX3YWZbt3sLJaJisTxM4XVN247MqYb+K
zNjkF2s3fQI6+cYir4BkyVx81C/H0Ajt5k+rQEIWmy3D9VX80yRD4JBR/lZpPyPulZElfLzHfqM9
t0EBOD7pqk8ff/jeF3w1w0+lVI4Yg7UbEnzeremEiEFv+HBS+pi4MOmGtvECN7l1ZhkWkyjpInmS
XxAtphe7cS1CcLhY4Gfj8AqdpctRsFfyfhqM53dXKj65SpbZv5iSmw4BXaPlpF7jvmzmvxVy787g
CKzX0WT0klsViF1cq2huXShvlQNeHloZ3PKYkaqTPHAQ2uDk7Lxwc9QR+X/u4tMncUcjShcgbt7+
KKb5XvGn6NG1Rek1uLhH+NN/bhBZgzIsqqLmlxIt119F+fteASo7c858lLBIbeZ7jo5NdVerIPcS
UciAJj6WqvDQ4rh/RgRQAWZy78NLFxCZH2ygpW69+0e4RWIX0/xcK5SwHk5PRQyROWlLDjC2CxM0
lBN9z/yWHPr4pEdSYTa3loX174VsPKXZD/0VTt1ViYQeLEc1lpVhpaOVqKoYCAAVUy+qrfWC5zEj
c+3+cJPTuDUOnMntZwRTrnJ+tAoZLfy8S3Px/UQBNeaJLsqE9xZAXqqiV8CyMI6qVjpnzfQcDgs0
9fezJDNOoXC9IW+iCLUWeiTPoCc/n7gqArEpIE3a6OawcZIRNHvaUcitFRQmVhJkIdpDAvwkKQU4
6iYcrANbj8JnUiPrvi8Iu4Jx+QGhI9Asmk0Z+/ecIZlaAewlgxkl42v+2zx6cnVH7Z0mbJiFEXGx
6Wv3tKawK7OmcOlUssZg7uCjjdiVorVoo1PFlP44tUGujAY5LTWCmvw8KaWNBNpljWcz5hDRcx4g
gDhLM9IDcAZy3Q6KaqMQzQaH2mv1DuQZGTcyK23e+8YwapHevt7akcSJTeflDNcnnxP7s0GeiP0c
ZwDQL+9Oz9n1yU55TzYINdde+fWcxXUzezEn9ffGFpbourRYamSAd1vhZPLkOhbQB5A2sdJz7Z1+
i0yzp1GYTPrMXoUSeZiHbGSRb6jTcPGb9Kri8HxiGwNCsMcnpgnZ5LmO783Mo56tzuQ01GW5isi2
Aue5TEmVjuP7YKO36VYEk7hO3rpVUtRMzfZB2JFzTNQhSsk9/vQMWu/vw5MyU4ozVQR6+w4ANhD4
Z5EpGYrzBWhAJurb+jrwRMW+EVbR5zbqbdoC2/5yf8P0ivnLkGcShJMmvQfpvdmDCgtWAZgOE7Ms
WTYVIiOY8/Atat4arWiMddsWoVyBu512P3vViV1hm5EkmzDceb0T+T5y4nuAVcKdlHvoo3AgZI4V
KuOgPtFJ/L6g3PyM922ZFUcuB7TSEN06XPpxRAkeTRE+W1+ZMUjuIMmvPLFYjm3pNmAimGW1zX8h
5RzITg1fb/fTSPfYZ+ZlkC3K+sjks8O3YVzmbMzcVASptNP2qYiJ505r2drIHYASMlr+P1bK+iYA
1jmjhFToo8P/OvGz+fPS3QHX3UQhRirUGZ9w62dAHpDNb09HfZXpwcWeDgSoHbGEdhJp1+8ayXiP
yPDNCdAAdHRmm6xHdPtT2/bsrN/g9u3xvbwWLf0XgTG+kQeiZJ8Z98aI5ZmYbEaZ5+JRBeFrIjc6
W8lVUpkSh0elcByndLz5HSbVS1SEmnrDdOgulJv/o81HOtbs1fcFprIGsnLiCK60LLUXNEr075jH
9HO/SYIfQv3OC2wmmS9D81NzQtdC78q24B5b6M5DY7fkzmtkZd9TWSU41F8fjrUW1SAZAOIlNwl2
7pTAVF1F1cIB2/nxY+r7t2zro5TVUvxdul+gcn7snXFel9eFfIXxLoLJGwzWQRdE4v1r48ys2ELm
PfErxxrWeUMN4PDUBerQd1ZJX9wEZUPG59EEVru8174qyVys4/NuB2w/ag7GL6f+5peOGr0x6MsX
4mKtoDQ4tqLZviDgvwtmfF3sId9x9Foe6YIFBoE9PCIEFduudqsDkDCL3rCbI3IYZbg6b0foQV/U
EST3VKrhMFiLI5WrvU5+Aj+AxLTnTuJcPri150on9ZegQav+LrF7C+OR3mc9dHrRS84lVVPvZY3t
EX9swEZUmNKBaKYxyh5ypxNqvYnpgJawig5jDnEK9fdNoRxQ42HpKJ3OEPbALS1wf3m+Cuv1SMaL
BCqFYmFcp8vXVGqIp+lJkbcDVWEjoQ9OHLlO5eZZ8fel6dTrnd+q6EbBEQd0C6LIw7p0dU1tS2lk
pVTMUfiYT8eIVgJz0cjjc6PxF9BhJpYvE9gvhT+tjd09fYhyO2rUHtTwsAu4luqkNMuo3Y0mU9fB
vdGLLldP2lmLtDHt1wifQQ0ZYRzR/6//boobKR3lCXjOxGRI1G1Cbm6Qw8uuIlmgKQ7wMNIB5XZG
jUDAlk1qvPSx76QlyqmJPSrjgoU9W88xVSroYd1ArSdxySS+09X34LOBsq+L8Ig/Lp/yO4rWWrin
Lv+YiErcy252UPwUpcCmy8ry3udUHFeC5KTtKdE5L1X7RNmed9Pfi8XLPLjOiUxSLwJ8LV489/Q6
TBlEHqgfGHo0Okfc+4u3MLnCXlhv9qK4D1MSC5Am5JJy6bJ6tuxtjFeVd/WGOLBCcpV1OG0PXdap
Hw9IZydtVl37D+egCLvl0lg1IDeRSPB8Rhuzv1Zdpx+4auJKrWjk5EFW72zQr4cTpAYLQpCrTQO0
pNvhcNuREnEs2LpiEi8qJcwPh195TVtf68T8/Us6f645zkBUeb2k0msadLlD39W5kYMB1R9dblMW
YIN8ZB2wSB7oddbN0Rt1a67RPxcvzkL61EF2NAt/DRZf0yib+l5CXmKYfhFkz5QIRxdtNHD/guxD
mRPqdM9/jdxqrZdjK+hmoj5syMqhuMvzQddIUyBXqDkU/cFuyV3I/vumdCDF7KhtCi+St0MmOkiO
/0bwAXczP9WJyRIyUklA/TkqNTGwwSlULMfSPBqqFOyaB6GwnxgxQKZQFchM345PeTC0jrfZClJs
Zyr+dxKUgRYk0mB2hZEu440v+E+YuBTqP9OZb5FtPAf5kKqJZGJJMMA0S1rI91eyzX30e8NpzVHN
/tH70ykJsJ7yZAeMwXXTSuthGXF6E99AY0gEt0kcAK/hIb8pJfqRs/F+eAeqxRIA/FIeRe4fd5+K
50i2iYRTCwiOquJ0VWhvdyWKPvgkVTi0iEWBq37ZOPNtAOVCtYZFsUzYE+6ZHpQSEhuCUzIzCaH4
RDA1o/OLmLtWaxI1qZs6DouNxMPw63Umvt7E+Yhvhrvx5aGPaalhhF8UkVFgMP7z9G2EY5jRvYWS
S4OZuuxCcDZ9TJp9yj7mBBVWSTA9DCGTUurwo802bfdEINBeVq4cghBM73waKM1cSNEOTVeeyF0Z
Y2/9mGUCPsMjL5qn7Nyutct+FltTDeVK6mpI8O82/rHdHHV4h1PVs79LHM/AETnOF7bzU//uGhwO
X7tAGKxU4UOC67zqCJwEDPE1ZMEE1V4DUn69D7PeW0nU3d8zKHbfWF0bz3e8CyNIh28hS8dVQigY
7dFuKEKwNPoGLnJ1NrGDDUdX6mlF/KjlXmAZKgSgIDxPz6yvNLsnWLWFZr49WHu3f1i61WsoeGpZ
fbXwzp+Fxm04gr9TAEYoyj0fESYRVIglW09uO5WZjy7RnNhqcuCoJPCmKdi4YEif5R7bU6o+63Gp
zbz1zMyfUu33BxNRVv0YfPKuqeKDDwLmhK65Dn+ZBUWetpzZMWcXiDRkONiZKqv3bARPNYh5Zbkk
YmZl33rSSOKWTP0AvI7DUjJ0iR6YCuhMz62DTNjgkNyKFfhj+YJ63rocmwxITdzj3COwycPcad0b
xKzPD4FDwzIY85VQXjzJs9sdfpolPuA9EAcyNriylpWUr2BlYP+VDGPHTLr1x53ttmSnG7B73ViR
EXNlPtNjopbwZBunAcVID75y87hk0Ay1k7m1N3GSl4xVUcFFm9KYEb4yyIbrVa2BDvMCJ3JwjPl7
DFXKwLMYCkItoYEAm6ufNrrOhQgeu2SZZEO2DIw3sI1w6YF6CZsnWfs9wtGEFeEvZu5ZRK30oMzu
6djaCKPzcuFLnSIWNF62AkPZnZ2pNeLVbXmUQnqYl91fqzQnGoa05RI46y3I53jLb7vPOb4/MRVM
dBb8TIuZJSilP6nQ7IVp2p8inpJVOYSTpyMtUDQTlX2+SMNfaIFBfm8/anK7VtVumh2tqCUxatco
MnjiRW49zL7Fq0Ug0DkYqXZu3DTI6G/AyoYlm7lgeeo2EtNnN5Ec6nN7miNAm4h7f7t3iCAJthJQ
e4xNfRxchNEuuj7SCU/ZK89Y+M8oXQxH2Qm3kdX1VMdggmPI0ZF+suegSj9Cx+S0dejvLp29eE+Q
n3eQ80rWTFcSybj9vxeVyZeq0zk683FIo1Ivc8PhxLANz9uBbuwUq+OvOQOMFbdutCuQr/7ajrR/
oMA4kJ5rTZPL86vXaCI9VYdOeYqwCW9BeDgiIHrMG4Pli0eheXAscnwI9uzgB5VMCCVzPPJaq2o2
Avdy7SchuNS3FijaUdtrHD62nsqWatODWJChC9RN6a+WEEKrwoDtjqmUg7me5NQZ/KFMy7vHDCwF
WhQOLZvkMMHpo+ZwJgMgLi30likmUG1ZfW3UJAWtH6Tjsslnvl3EYOKgQQhWW00LXELAYQYjAA/i
Du9gkl2mLwmaJr3eqqZr7qMOOVB3g5enFkz03I7CaWzdAAjsaQVBNrIb1+CLU9sAxahEJKdTfrrb
3NWYvPnsgKmJyS5MKoc1QhSXKx2RgKx8ajdZQ/bWuaKAH4rHKYSRwmZ9QlzF1yFHB044+bg6eqw0
n0beqakmvdrG4yndwlssIlrwDfi8jfNuZlBC67NTrpehe6NZjuxjWZHBbXHJTIFQyA+/vmVd6lLu
OdgkNrVxu+hgiEburme/P9UDvEbUIuZ/iBIIv1hJFzbkuA3WUOSxQE9GjkMEVTPa8HjVX4tL25QL
OaxGYXZzfwDamuV4IF9Q26SHbhoHUd98Q52k+R/4Ay8ynbiMZ3Bdxn4dmx8gPs+pFCOtwEK6W1yA
OqkdcXRSF6tl1i4gdrhYtZE0L9X5xI34nebAs0WtvJYqzFnAgZ2BEXMGyD4ElQvR1t+Cx7hDms/R
xAUrmcyqcR8ML0Yper1WXtgGsWOqAhxfSwnujVVL6rbZ6TTOSGMikUb4k3iURoY6IWI5b0TTPEb6
VsLplOtN0z/sF+nqLWOI/Ic9BR+1KVSIcBQafiiARFeL7g4LIgrwO+6dP+u4M8/5IteNQ2wk8sIH
NoyZfOAEUaQfw9A4apdjro8WnUKx/c/q4sp+RDTGziTTqLGfwUWZPoYHfQr9/xIuDhTOun5fpgu0
jEMLwSvYno4zDvBVOcuaLGwKdKwnZEDSsMzpCFnvEFPuotJ/0nZ0Y/rcwb/meCMd+d5DEwu1ZKol
7uEY/JSzj9vriI3n0Kx4rIKoi7CFtBOJEKSIro5uM2j/Jiu3PZcCraJlpzyk77MuPRcEGz76yd/r
dwwA+2NSJZJrzf1x5vxwptw77zGWL+K+7unsPSVEin6i9fhOLXyden+XwqZzmTowXDFmDdpZq4/0
MtfxcoUAYe0WXEl3Z/4G3gEZ8kGP6dY/yu2z+Vv/vydreMFrBAqVO32pMUq1U37PRlbkVJiGyOvn
Kkkc9IagZHRKel+efz7DsfEDrSovfu9govBaCH18QeelPK67bxY0QWdCdds94uvZk7EBc8w7zw91
gum9u9cUa+cVKf27Ne1RyHiiaP+03d7ZOTU1w3wKcg//JOTtLNjnBOfhFEmtrI5g8X8KQjEzIx11
q4bquScpEgy4IehIC/xc7vqDsGF5bWDBT5Ey/ZTC17Dv647hLRJMn9XTmsP1OuuBE/FTwqUoynYg
5a8O0u+lbkljIH+YDBP6JVT/LYp5ocw3tV+qB03fJJw6MNp3dNptzuoaywr+l1YBEnYcsCXMfZfJ
7OKGd0gvX/5f4nLPnvOAQq30COA7jfhv2rOAznigSDa94FeWXhM97aCnoEMpS7cwuLI/cbxFJKNM
Xs8+WF8iMlpx8mGYa5Jp67wDFQiqCD+ObNvxwqGTudIHY8KHzh9AKEXHAs/vbUVdjtkdDoTq/d5G
NyaztgpAFWl1EvTNztFmTsVpngc3SNa7kmyYumh1RNxu+I+96rdrurljOKx9eM4Sbyd8GapjbFrT
LXKHiO5smkky+FxRAW0+70N+sXgV0mCXOmtG+Pn1dNrNO/+aOt4f/XlKqzguhvNw2zo/fdVqfZbu
SuII3+JcIudK2zQ4lG1EGLpF9KVM7feGJj898tjIQNR0hrKVAJELtLUpNdbATotGU5dbCFJs8Q1V
m+H97NoVgdmartXUpJ7tP/WBWvMq64atyH/cy/621vdOxTSpVtbAXKwwETgHCCOA3sFcbiymn2Ra
gIyJLqPaUnfDRQfVdCOmByQBg9xk19hxlIQINPb4QcjCNMZ+m1OPGcwiishjHWV185+56EDmund1
Le/CgoccrAIklvW2DI0B2DmOroxDQ03lS+kdrF+yqACl1dIvnc4rLRaaRAQScs6bICDVW6ef721i
5z2cE4iMGoixVb/imGTSlWTkU7CECA/Yrb/SS+2ZTZsizZEb7uFWqS8SmkRV/rABa7YhHP7vsx0Y
jaInedKo7Kd+HNekZPmMgp+4ehxRTnbQfUCuoTzj5aEA0eVX4PKuvBsym0WcTpZ8Vt/zsMuX0nBc
jz2rJcnqyWrmYvXswkxy2NKD2YCkiJjRQG03/D1eJDLcX3Yd/ujdCVmhWOtoHeAASj6ISMgWKXmd
Pabm09qUDlJutNUW5DzCNk5xxxjAGPxrABRj6rFsChT347safxabfoRwXyx2OiGXlpFai4AWjDZP
J1CAkXBJFMhoaqDTPlRB4oJFu1L2q067KA/l2wQtvHSqSnkYH39maJMmMLpxanlDU6+75a1MNWM8
gst2auxJXWrMFzCsFaChmDdTUiuci6iEPBpX1T6KkbXN21hS3BrLR0v7qLigB7VuSBkXyFxa1HYq
rPGt8rVa07jchhC3RTIrhs/tB22O4IMHissTNh7InCJu0/UkmWboJhymTJ1peZfqptah9uC6TDdG
8AZjPPWoZaB6VGSn6dJh1Lje6LbEnP4rassbp7pfUISDpvpxTCsiZPrQXQkutby3z1A+sWmhBJPV
skGdJOvs2AqKsNmOKql0XSCc2zzXzr2zRZ2MOz8dYUTXsrGCbJ772i17j+uGjkRAW96U3imo7Ti+
HWgNep4mXug2LkwhJD1+Jpo5hvxFOPZouJUnpROB4MFBfWMWsIMu1QdE8ILNVtw7uysTdVkC/HtQ
kHaixy9DNtMKPGG9Far2rAfJcySAkyN0Pf2qZASy6trcaarbDKDkZatMvWoy0epq+MXfxJMhhRGX
JDDOWOsoqhJPlJhnYH3Fvbdh2R8NIrQnuDlKtM32iJdJ2Us+JzlGNx4sSEChopYaiGp5m56l81sj
BiBQ46kL8nrWxNCPdOUfhFhaVKnjOgMucVkIyyEFANgEgrXR+t21JOiub+4UdvHJ0by64H7RiQbC
U0AG9pBVtYfHCKLRURy9WMwpwzqYI8HvBeM8s36DSTx2V4A+CuWL9Vb2B6cAD1z20zGWBRZRVfI2
oWr/88pkfVTonZtubGNw5NTc8PJCvovfGm5t1Vmnt3pGnAUnb6v8HyFhhDAai8roTV+t1XBdycLv
0+faFkTV/C11wPu/XarTizm29sgpqkAWGrbel5gPRl2UyjaUbUB0laDAmZEeflWKCq78D3Px+G3F
qWp/cO6ow7/nVdueUNUEB3/BgF+ogVBIvAM7R9P8Xvq3EAhXM+CS86daAkqz5XQoj66SsRBHZpeZ
F+rvuV/3e114rwkcQsx8bdwbiWaFY15AxK52kzEYNL+ISrD9ogFHe1lKfexJwECHH5FLC0T3HGiH
lk0a+12asNsyKiPsRO/YnJNezByOGFP9OZFUzmHhqVML53feuD5JvahL1c4HScM3jGhIiJWOjQ61
7w7cIAolTaR6bcOtDSTl3cV6oIiC5SxOph0Z7rXymN7eouH7XlaeZwiYFC/Or5H49Ut2K05Mtl8o
9ljtvLBgScGQbghRplWVbnw24BN4RuTbwmp3F+K6QmzddLPRQ8ObXZ9pfnju/jGSpjEpJfJ4WNKt
a3nR6kCvkKN67VmFXzSUWXDXxKpwy9blfn+ozBdVuf2lXxTJaoUj7pGmpg9QOaxSPEicHkFh+ZWc
A1TySN4EEfYYdLRD2ooZgsivTqGaBW28ayMv5Qvx6eKWVcp651HsMAaGRdpCAc+w1sia6+7V0yZR
NMS3fBzDDMjtawS7oiIU01IpwZtflU1l1XtvcxRtUfI+eua4HEfFrqYkeSTvs9EBdCZL+XcIv9IZ
ofeW8UGouFPeG6pyAFyWmNvrRsY1PzMR5P43YJyklw+7KDCn1Q6futI2Pi4muhKUNv9dAUu7u7vT
mPDYxekSp/m8ULr0QnxJbT6ph4iH62/HENFscGfyHAWDnZ59jq1YK/otGDhWqZ0BCYri2gMEK9uz
xPERjnLRlx//7YkboT32kriDd25utpNgjvhfyep1+jgHkt1+b+2TfF6Cu4fPzJz37Zni87+HsMWX
utFUuOjUer1BmMX4TNK03BfnkzZY7Lx2L6zZz/L5PUJRdzQn9kC7jS4409zt2lLz0DVTY+JWv0py
XfvTx4BY/M5gYTlccJ+PRYxVevhCLBj9ZmzAJQW/FHOMq5CpAfJ9ZH8nwe+QMWptwkYRk3q8dln0
FBozgoFlhoALBW7ENr1AWTF9Q5z5pYwIdTc0q/mx3bum/Vpy6DoFmibcSZabJ7Gl2cdB90sixw4l
nLG7DvRsEzKNt3N9AnpBXFrMdsFu6B3mZok3kOGTn7CB84FQkjCCFqkMroh8yw0Jh09+YkHREx8N
fd2zit4dBQx3yAHQ57QpSmAlup6wPnuSyDFKAbjehkLI9gUSsHUUDKYgCzeL98hPX8vetKl4h6ys
3z+whtvb9NmWleNLOpBQ/tdQ7AZp4jhsINgAEJ+sdPyXz76UnlfljXFiF8tXZoUMRZg9aeW+b+X9
s7nDkhjxxwfrWkARRoSDuhti3N2adQNRs8d7g0JBBkAlrC6VKHr0gcmGuqe3oDwyCObmrRpJw1r1
3Pj03OME276kqyG9glsiZ/9AP/WXeoOKCujXDYFBj/YbS7c2pGgl6ENEXSfe+jsYbmNKF3/s1TZc
kzQol2DqEjLVbsX0OLocdFaGrEd9Wbquvh4F5VkOIexmdF+eLO36VVr7DLHZ95qSQ0bK/e/18HrB
ODZQg1ajJX4Vlupq6BfWEgazR0FoTxVVnvwSqzSHp7N4hAuv8r8OIIro6coXHLKqtJRnjk8I62Fl
pnWPbef80Pq0cn/Xm2sZWEGjWHsjELhbGlm6xEUfHAtNsa5qbjBcda2MQOcu0f8ocAWPs6uzRHJl
JmkxIeUqx9nB4huz9i2+I7fHevLhcbLdGt9Cx7KbKj+qJy+vi+Xf/tRtno7uLJ8X660HF5dDJSc8
65ZK/uubx/wpZvMRIN2epVO19nHya6SXy/eRPAmHujEbiL39HMGdF5p6+8hkIYGulhm155EoUT/F
KsIeHxBDcf0QcEj3lAAaRtVSAhK0zcs2u1RhSzm2guBoyAbCG+05+ScjmIO7uiXAZ5sstETsKxnh
r3RxAaMuUTZpZwdymUKJCdDUwaojBOI65pqC4+BDCLIULDqmIhHilsAijowIjzNAB0uE1gxG3uy5
UIv1lULmvY6108zdWE5CuglviM9PUpgzHhsbtOfnBM7VwvwkErNEhcGuk9efVAWsgw7AFTNCJ3bd
cR8YmcaHipqdjBbAMKE4rOhsBBHaummFN+dKZIPS6gM9Z1w3g//DG1wLMMO6hZYGXM7703xiAZpv
A/ctB2YHqo2l7fGqwDBg5M/qgSuxH4jxqlRl/ldyLfHR8h+cAIBsA46hnWwuzZ998zBWYES8ujmb
8KXMztIoS5mEFDvT1X3nqc89T8RDv8RdSM8aewaxWScoCu7jtiR9JP7gbu2RwbYBom4FDAk2/UMw
YLmQRxuBfkPR4IMN0CbtGRdHlGJs2aMIUBFUXliZIfZazMEKXwwG6KC0d0aQw8ZfdY4oZC7uRdUe
IDjUgoR9eH+msfq+WaC6/GX80enSzIEitN/yLJy9VyfKW20lv7+eQ0YGz5ZVJS/nCfCwltwWMyHI
KiDmde3uD4uP9m3eyy5gWd9ZoRMctNEKFXPMu/vLtV1b26/FYVd8O8ZbTw85XSkEWyDNWsqJvBTU
3yqL+I/hHDiswCFVIscJAx25WRdcAFrj2SyIo/Qxy+gWg22XKkUXBL3XlV3ItqsVzdlZ8cK+AH2D
YczCl4YYGece8dAJM5FxfCOzgHLjRtjCDGPAaZqpxZ9MiQRPeNJ6MyCvv+tkubcakOlQcnPzoGqD
mSvviyQtOywM8cvTx8tsFDV3HQnNXziLt/O7FP2V972eaGBqCtKLjG5047X3vnpG5/wQhcTy1BIP
aSzRDatez9qZsn1MZRDcBkSDfxm2Al1uAN9Mv626qjAlR8RB7H+KReX7BjnbAzvMoe38ZbKRgVh5
Yoeli9izJpPverqSIO2ranhWTodado17qCQVeL3Xx8Z566mQ4bavKR12+WK9lEfXmeie2/InhjzK
akzQCAj7+NXqIW6XWEfRpTbzF8ksotjJ6Y6++D8HOjvvZh0AF6PLhMQxRYjzNbjAUl5PgP1ho4Iw
eR/xNfgN8pMNRT8owgM7g3hGIWxSJl/F4pmxDksTIF8eFQd980qdauQy01u6etCFY8fZ6rqb5kXc
VNe9CPeMkJfMtyu2Jm2ArRPV7szAyzvwlCvzmj/Uhv1RLB9fgkWNEfOWdR/WB90R/vGuZhza8Qxm
4wBRUnIwcyyoHRhCvo2lOJfA/Z+X8O6UfrmNvaVwkevs0ykMoVsrIbIbJjCAtxF99d5nphQ0dJZC
FWBFybKNXL8dwJMu2rPdW0ywnkPs69DSEBObZ04DNzKar1K9wjya020yoOc7/assxScr8md5NNwD
Btxk/H72HRfnj3C9W4F6EaSPzLCW5O3VaYBYQaGsVHw/sM5OF0mRQRM6473J0fMtgDOwxIDEMj3w
QaZ8ureQEAoftWkRQwA2nd4j5OlhN5sWdpHpW9zksEBtZGLYMFGYCwYXIQwjreVJr4WW7YJphUmm
WgcMQ0PUPCZm6YuZhPaysFZy9wNgn1ymXQF7PKHH/yp+0on1qpkahlNfHrzbaMxSuDo01p/cZrLk
2zIsSEaUYEllcM6XtlEIbaJC6Kz+xMre3qiv82cAwiZP0kQkasc9tFhduWijwcOrqT0q9hWaVKy2
uoGspqN68NqHrY8apjFsjCGaWyfDGu34YbIkZHzK1QFuUmwPSewsjooRP1QaPznWYRd3jXInRQGI
X3ex/t5ExyeBzAjNsPz3OKvS5kTgLi6+4NczzR3Uf9W37GPynyLGCr2nPrskAkOyDX+5sfRBcD5o
j05apNPfySbjHNMm4It9oVEy2Rq2TzRvvV+iJkXUN5U8Ag94zUBiq3jC2dRe9R6ZqJaJWAZ43mgv
2CzVD9Cj+ff484PPF5zUCgn+o7sf89YeuRe1f/WOdpxK8TpVTaRXRZDMPNsZCc5JUNCIPPAlTn74
Hz2rdSvdLk9WvCtFf6QGUMTgDTK4ZL3aVSAI5Qsx0rKnjXi4Rs8nlSmSl3u70pE8iLJqP/W9s9ke
DsoHiXNpfOmz8M6JzCXwKc1R6WIadgQ3UYtdJXvVzNx+7V22faT2Cx6ZXxZO8Y1yzb9rCQui994y
16DvurvZsCYcHx2vJE/15Sa57xbd/d1rvXNq+BvqRWY49kNHbUd+BlhNEaraMG2C9gnZlFZh79c/
LoWNgvUlWfJDqQ+9ZB+ga+jySan0yzsbnNzPBDWRQ9SPa1TnReDqdWsav6B6hbvQpxFyGwMvLxYh
ETxARX1K6qWHyAgGpsCnP7FznNOI82hYi5349vd4JrdaeoEkXIkA5/XRPvECdOUs7f6jvXuPX1Rl
lQYRdBPSeHmgct9LdZbJEUzHRhvMK7mNYlf8i+koA8kDmhPAuNOkAggH+duQT5NcdIneZvGhwX3O
2lyG0qZUnJWPiHOsUsyIKgoxLQ9mEW1HeaQZTMgJTxDxyoQajapVhoI/KLpMhrmrJclqmZOcDj30
I+SdcNI6YrUTkLrJgiBEi6Nv0XVvJVAzyrnVW73g49txDyXKshhub/t6l2vlecTsSXweCckIpVkd
NvpDr4S77Nlm2LMUV2j1YywJVOw2FClHv6poG8A9HxUuUEeVZWbkocM1cj5DqzE4aKdl5gI/Smua
ixmJwGGGV9eKOaykiRwq0dhIkqLpEBVVWTkow8Eb/t9ggtF3Kd8M6L7/awGNDadrH+f375G4b4H9
Z81GPbvqGifFN5tc1oZ96HsZORD3pX+ln9AUu/LtF5fS4srNtrmmEHR3H0U0lTK1VmLmEOvjchMJ
kUTqm+MaTtGYAaPEzdmsrdYSKjY5Xt1/bOUrGGXvKx/coeH1onJRjCF3Y/w4b+Y1alWfY4k3aSrg
ySLFDCXj5a4DNrofQZtrli7XbYex0om3veMuD+WKW4E5PL86lNSR3KItJ9niLyebGRXo0AKefboY
6A56Qy0nw5CPXLl6bXjiJ8nuQiRFpcFBaaUZS+ES2U6tdqorI/hVQmXavYMSiGF57tUey4CnKE3v
j9E5jpCOXK7hQPerRpmJ6tULr4NiiQtyHIjLOhawMCshk/rcYPB7FnguEizjOmmPaOUxfJOWLFrj
zHwz5z/jl1MoCR/jDgUgOQhoNsooEFUmw8zbJSeCDtNJqctoqu91pRHX2rhLfuOAYKMaPBIWuC9k
4JOuOOYGB3yZqHl/tj5mSCvOr8owkmHWwLtvRLJoqe29UYZg8ZJW1OzQ0RzD8+0Sjk8Xnb2aVAiE
5SG+9UzULMqln2NBQu6naPac2aTvKifO4+AOcaddvnB33ojz5bdH75tYqaknL1KJTge4BqmtEGye
KNo2catyom6j4W6l9jugt38VVeDeTI5xI48WTc8TqrabowuqhtQndBhfBfn7vcLILEeP7x6XJGcJ
8esK1S4EkGAJ/DNw3fuS3Rw9z4NZ4xKqXIehMjtYLIvjYCDrGA4nGDsXjVQDhIXf8Xo8Swzt713v
XeSyJ0T+hpgSMQFY7C6d2fmOcnyQZeOD1IW0MiT4VqgRyBEWzSwqK+EC/bgmY2ICAd6wTUHI6/X5
eFD4yCBxs/yNIShMSEqvAEGFsn/jrWYlp9FyHpQSeQM1HUjDcGdvD5b+qTQsvuqwIFPMpZ1ixB8/
cQsiZiqXz9FICXLl5hlnOdd4ZsGOGJZOBxuin3oeUnJI7DBE8rOCcsTlaUV8SXpmDXL1DIuUGSIE
lkXTf36k8EbEVzkGs89UKlA8lE+wYNMuCuxBH/nxUpfMPKlh7G5kkSxUACl5uGKf7rwFYpdQAFX/
hbIuPxEJ9J4cFEqjq1csJkH7JLDYLHrc2mObVYFqiSnvkL7GAy03wmJCwZOEm1vyYZUnG4hrUgOl
NRzEzR4IO2VsGuknHSohboB0/rFCVfigog9R9rtTSpsm0GYNK+LAApcKrGGAAbTcxL/3FPbXj8jE
BYGmoV9MLYAlfA2h1cnbXeqhnRvmXruSq9nQBG4rSsbq0IgmAKq/U6nx8iSvWwzn0vEhTdu//16X
02MlZj2i44sawzIK3V9U4PXHiNbwg8NuVFpHjScxT1OVpIvV4AvZNBN12Xb8vdLcX7AIKec9nHBB
SGvo4XnlctFOOa0FmgcYA6nOV8oO0e0neeFxT4DFtdYTdBZ5pZYmYZxzA1YTOqisbWTzcMGMAfs/
/WktEbCyELd5st6bMJ9girTdTx/B76nLwl0mYcOmbCSdIsFs4mOEajOvzmbipX4G+D6Q64/PoCtI
Bu2Eyucq1AdACZHeyMZWlKCw25dyFoDlaCG2S2ceMgWLVCPeywNk7cUDUb8EON07sdSuNcX8p15/
lgyroqZd081Fn6IXUpEJA1ZZeiU4qmeqAhY9L0op+VnJTjYOLai1102brJIwNpuj6U2nPEBS1JYe
cy42L37OIBYt4eNRz5BYbyf2i+oODE/Vh//JDOwISYhKgiymfEggsGcpGGf1QwxgAaQR/zxbp3as
0q/saSYRyfpy09plGAUABg2SsjtFVOlVfcGSSmmTZnvCFHg0705KC9wADSa0mViZtNTztQDG+VD9
9yBdakRpvOzLlzf4VltPTEJuWYWJUYRH3tdhmD8PwbxyH/2ga4uplHCT37zHvb0pIsy18jPPHqCl
LvEfq0J1VHqtJYrTlmnoqc84c0jsYKq21XihEcRpoEZDdbc24eGnMsADxStBYI1ecuQ579lF1UHA
vaN1HmjVLjoYU3mV3Jvq6Dij37NGYfP9Ns0RyOXtoeSaP9Bb5dXR2dpsnwBr/B/z7wuvCbwKGEBA
cVwRschfXTgJiYVAyt5cpl8aNZeLJr3A6woKRkf1laLWn/LyBHzL8unOGDX7esJUeVOn0aJzCDKm
Q4unZBujAQl0/0YFGuGQad1KkJdEOrjZ6HYsVMQ3zYKGluPjLdAcEKrGy+gnVHUK+B+o3lnTMrkJ
50so7fLZwFbOEJtqG8xAF5YyyulEHZxsWoQjAa9HWwrJONBjXDzi3y0FHQ7DTt+J4kMag5Xj2Hj9
lRd5NB6kzZl8IULxor96MIneHU1LkZuj0p36CcjGX8xpX34GaNUKwtToT6kgvJZfNW/orV9rQ1Hv
FtLVBZjqOJuVjRvNNgZCMEdKgO9938kKYdCuJ0OkT79nbsFbNXeBsfc4Nf6E6c4re2HDNXbG0uJ4
F1NhRyCWnjRlfbSEsHBfI0zSUNbTPlcbYyVc56g27CPmW/oF5tHdIjR6SPJcEyNwDZqT13m77FZI
frFM6Ajl78SmFd2FWLACFlzMKbBgr85VwG7hDwKcKbjXmxqe0oe53F2nTxLsH09xsQN8ZELiQNd7
cpTQ1dz/Aw4QuJuqJBkhk4pT00FsdHPSQcioOkHqoibeTO7ZTkyhsSgZ0/+H3mua56nklpvRRKPF
dcF79yX5iPv/KH85acfW1NwAW2E5hqXwmzm73PZIIHjmME+TR+xtfiaJAv4qU672fL4OVqsGDt/q
1BYdVHIFIclbr4O1PdLJl7W5rVo8AK2E3OV1ZlaN3MhgeXAASPb6knCHoRc1KorYtDkcENSy46VG
IhZGZBTtVKev0cO4S7kaWUYPHZfZjNSX28mcgXKkdS1EJ6wruxGDtilwPNDiEAAGc7+9QuxnUckC
LppsvCh5T81dkOnf3KCxYE1Z+nDM/sq/sYPlVwGud7CkIRk3+lje7ZRHVoM8JbHoVHTXdkbcJFqx
okacjlZIJsySoF/OY2CVkV/r+DiAXdUmby86gDuFwadV2N4YhkBw1oocbSo+RjLpF+iH8ZDajHU2
3lEgFgLOYmOigoqM1JxhfG+fxQU42dF7lYDvaSSFuhhZ1bed8tzj0oqFNRU9qgm6GUwm9lX055oX
MDiXgth/UYXfysjQ8kEh1oJjHZysyTUFZYqis931D79yJjArQKKbUeVOYfDwsQG5sY61A+Y8w9S1
9NQINaOyrAb3KWZz4fkMlimdTQVbP11bnBlSUYuo/fV14zBrVkBKPWUU3mYFDp15qD9LpcXvFAAu
3FeyZtXkjAvVu4njMtzkBnE/AumEPsvFUT02I5tawtCOPgFHckZ6KpZdzc8IR5xpIzTyEzY/dKMK
vNNS4sGPXPLzrRBt39ui3fKY8LYC/pRmqe83aU7OfaDySyFDe8FnI/A62vJaKPjHOrz9Mzb3yY9K
dj5d0bkBThpD29NSofXtvOfjy8q4yXSAOe8166l4Mpx1AEZ0aCMDtpFN7zDe4pEqhA5RBZ0IIeQz
79thYorrLkQhitmGMB7YGJtBek6fk40aukuhqz+J+jGvzwH5V7herupG9OU17lgvunY9amsawG0G
B23DNcbkSKbZfAL1aqPzEa/9M9EFqSAEVg7/RyGZekX3696iFmOrpG8q+0XGlqVwc9PotC4yFnZf
ZOGXQ72q9RYHHzCoMdr+wlAsuUAhBWCnnXIzizKcDsuaoeAbbdDzf/iKreUWC6u2PfMUTPEDLwp1
6HDnxNpBV8ALJByTmnGy/+wJ7mOg33wtifxNeKKGVqX4NTg/VjsORPxaXbUYX9mHcOpT1xHzuELf
iOJRecjKDR87w+/jTBaYTL12gmG+aN+sfvonDd30Kl10uJv695P42a7mhEvFlCU1Mchgi/ahpy4N
0Hn+s8gBD7U2a3qC9jxhQvl7VaTeVe44rnky9VQsopsVUlUFG1JUX8wT/V97gYdL+icX5JIlDUog
l8HkM7uolftKQ/gnj7oM1Gr21qcp45RAueU/8YA4HVWoNeIpwLe49UGeRIxSzHpzp3Fh6cXQSuZF
ehH2U3DCgYkOj0KtVzd6MlqLk6lHC6bh/3Fy6yXoNUI8Po82dFTEmBo2MVd3FjImYyV4IUGU17kr
PK7bcA2s8o9qBLowZmffXGstP/KgYi1Z9bxsRpkr+Lfhz8zqzy01/J75Zil390r2dDWABZY1z68j
g6Tz0megIie4bcEkuQoFlvKswHVn+dfF/eg3KIZupYrJ+JDesjuVLrAV661mA6b37v+BFqWo9iOh
4y2wso8jwxNAQMcJLMvUVpcD7QEOHLhP/+nuFvmNNG7UKtaw9i0eunI0OEvkJonzvDUP8ZyIkjnJ
FB8HRow/oAzw+Ih8i97L+FeUdGJon2BHkosfV2YLWGZaJwVSGxZG/c6u9ITYgvlRcdvZe0Qw7idE
2p5a5FPL8Cfs5ByOxoxoJAVVVET81XOMrQ9kea9e0kqQJlqYEYrL4G2qxwHdLMRoA/vfbcG1Zj+Y
vGl040Ezpm/G0lFfINTcl0ijTstS1/DOD6U94sHa/r8pqk+LRn/aEEjVnWhL7AZk7f7FQAQX/Q4y
gFTJFgQRKNcvQJo56r9OswWhak64FkW2Xc6SkQvBztU/FbDq7DtgUA1RO502nlO7Dlpnrx+aNHuI
ZijTZEJ6OwnUv9WrKZf0BiBM0Sn3z3H9uM3LvWeu5w9jR9DcpoH++cP31Wzx91I84lVupKP6GBk6
lVX2sZwg62JHIIv891Mx3mtz2a5PYp7YNqPxdUsGjx7CCY1L0qpt78EJN0FDw8WBfrClY/L2A8g/
l0JXWir/a5u5imEaUGwQB9GDg8BWIw0lkV5aL1DzJJtqXdxBPG/bSech8spu47P2HIzd8sgbIh9n
zKuQx0+GQmwJBVbkMHURlbsUaa3W38ZIRjC6og2uDK6PKCVRVBEsvLiwgyP/c9OD+EN3BaFdcrpD
2aoYblZUrMfjXkLjxmh3EPyM17wiLcy1yE+qxlHh2d+5ML1rU2UHzEPTdgaGRbNGt0hPItn/xNZY
9CwUjlGbU5o0TvdwytaQOkasHxMOQjdUs3oIMzZOVELO3AaQlWkkaTL2ALMoMdUyZzgkUDWwCz8R
jZ1EW/QZfRZF2PQAXtELLDuQm2TiRo0bFk68TAUsolROcnLgm4TZwxHFiFs97BswX+VhOgQcvgOR
Y7VB1xpY63VmMKJ+54Pw39VuYI3S/UPtvfPEug2jl34KY02M/n7c35mfGmp4Rgs45Odn90W26T28
EnOeFc9uNcNNl3GPzPomwHqNz3bebp1i80aTzaCw/KXOt6BnBEvTbdYQKX4pExOOqXiXFbQaWmbo
tn6Zzo2VDEyxr/9sitP/onH3zqqFXkoT4N7HjZMQEab5lvYyGfabMh6NnBOAZHCLVOd8nF+8DtNZ
YUOR4U83ZcmqWrFxadVREUiaAkPeAVwERYu86BpvCgqupGDmSPyLV2TukmIErcKgTBkxoY+2HGdF
M+2z0+9taLjkyZ7qE4ilzRfOpWS3F19t/KdQLW8ivEz9hk62xfRUXn7eH/u2XxX14hyC8tFKrdyh
HlX3bDTljGMw2mnOKLKvWMXL8jcVCE4SyWJmg+/SJXFmPzLC2Lqyixjh0s0yIsxywdY5RGsEHj4G
eAGHuYnFq6RPIEb7ZJWkGsrzmmGRMC/Xp5Rxc+iWHdMe4d8SFOfAbfowA7fDQqy5MeFADuMb6FlE
TE3seBeQjgi2x4/voYyTxfBUHI5wvGG5DzBYccBz2oebig/pZPpkaXAxr2f0vin+KCv27tGsv+dM
kB93MCzRG44oXlVcmUb2eTy4JG9uhDysJl9msdsBwnt4lgDWg39i4FaIhzrAjpNBG1WHZFU97UGl
1eGxSNNrOjzvBNorlDbEcoGNZNwg2e+zfZI/4J0HOViNNDytin5BcXGfvBJUhfwa1LvbSabOUeZ9
a8SENkBFpWlk/siOcYFq48APUCu6d7/L8Ac+F5gSARd8oGjrmEvomV3aUDE+XMonNLUZZYlvce5R
M9EWBjfKsPei+8bKexL2AwQi0HrIBo79Hitvk/S6F8cRHuL0XVyvJ5xpHeIsvJL4dNmiLRsSyEgh
DCK0cNartIPRkzU4p3uFA78QQnoo9ebboV1qGFQlKnLejiQQHRTcsDAmBiUuvvCOYBFC0UVHvOzF
VZd9iPAj4lKG8HXMTcfKF1gi03Xs4QU/5PYYUW4sOgJgBVce9MBy94wgGPXeAiyXnhyhMw6fs/3n
Zs7XB+IuFhPwfvDQDJAXZE9M2jLSGIVhGUpMnaUo3IiHcY9rvAVKZt4LmM6qjpZb5Qho2+JXFlI6
ffHvFWN1YRt8wyX9n7KN+7NdOC+13zvELwbA0ai9MRUfYqogn/Z6OebdtmI/4EFLYNuG5v7F1d8i
w5eMtWuSh75/jjNbfra+SWxvZ0WWMPtKmi67i+eaWkmlxE66RS29Oo2ZOGB7sKnyhKePj5nvHaSz
nmpsju3Pt8H+TsQYNkIEmbRWLsuLibtq3Ckb1jH7256Z/ndo0kGP1pyc9WFkQienldowydcv8Z1H
kwgiTl36AFDwZ7puQ0Ua48dTm/oSYxNcq0lpT8sbaKzn4kzlv2gw2e+xDS9yh2nOVZu4FlSEU+tW
ieR4jNW90xGYVOxwbSsN/sfonzb+0T11yPLWg4FLKdQiTvz2g+Wt+kTmA5Ruia/oI7AANCMHZfWF
ykdXrGCb3u8taQTHMI5y89gHra9hX7aOLkUZKojOR8QYREhcZjlJ8IkKFwR1SP26JkV6JuEr74uc
JeEilh6OY9L5M42x9IKLiXQFlbQgoiRlysK1GO5uguzlQjoi5sFPUkI4HG5pHuZJnv8zPrHFuaa1
d4yinI/qI+aFpIa9OO0GNoK/Cqc0v/vwI8GoN8gfReW/0pcbZ9UVyrCI5+gM4Qaq2vGvA1JY27AJ
ZddWKhV7irbsBsh8LOXS8hX+/+dmX0DYd5lGW06rtywGg322yX5EzeIeaGqfvinw0/jMUWFhy2bW
iuC6mtIJPdpA5Abwt7jmDVkkpanM4c4M+3aMsfSHZqrxxZWBPY7Dv+undcMSCaJAhJ9619b5Iksd
yXN3n+BZBZzS6NsMknkbGnyGo6SKS54G714FDaVIqclGWgoJ5wqhqilAZYU5wKuqROoWY8f6L50L
wiWfH8AdLVpPytYlMlJYCr8+ZOK5JKTyFEsyyFlsKa7QGsvAvrfkh4r2MIZ68EW4VFYaI1ambxJt
2vM/lv3Ls3uc5z219EuT6cpD+wKMtNW7sjRsvh4CEkMj77Hhno2tgArIPiiZYBh1vfsS0uzZTzD5
Ib7rsEXpdK2PjXYiZWwX1w4jWnVoXkcxn93tytg7OkbtMdSgzzVWEQVIEtW1SS66oKMVVGm5Gs/c
9QaH9xNlHKEghS8V4WJPgoMtiDSo+wX/OYneHrQ8+MU3yET4dXfbqLcqSCtH9NN35TEQfWxF6qvd
2gyYhceHhaVgxuZZueq8IObE9fcvd9cktlfYQh51dyqwgtXSdHIr2Xp81XFZJ1QZffIqx4YD9mT+
iDWjiopyZyqvEl/h/QShgCocEVkjhbcXqX+GSdKO28IQ9ti3/EduoXXJArkgQYMLGteq2LeEyTD5
AkUZP4ZsHdIhGxxwj+uxZjInNSbgNEdPHmAdg294WqcmWRXh6P5QNEsrPtYEPT/EjZ1LdyobXMsZ
H3j75srKeuIb6KK2L4y/DCrdz9XpOMAP4hT5dEoTAhWO+KIhfa7zCuoL80XIcVV2JWX3DKvgoHNI
q9gYpybjqAjK2Li5jC1mtk45HzC4Z4GcY4Kso2MFqjPiMeQBRCppXWZq2ajz4kXpQnswwlhVJavC
bZSwWuZclaQ2yWs9Pxx6pRBzDBGMoF7PS9rZJgMN0bM9i/9YfR5gc1UbMKkKensZ9tc4ZQvwUpJ/
GZvDJSggstEXk5ICvQfuFbt5iQdmR6cSK5vForm4Ll/iovOkPdtp0uBkVxgKn13S2MhioJIR5fD9
Paz8uIgFFeny3DW0uq0nqNOibSfp5VzGsWLGjJGLNSsliFO99Y7Ze1a/YlUVktS1myv4P39TJj4z
9r8i2Z2rQgo2V+/CKJNrUVGST81yLkSO6tcbsgAHeHjIwiYcfEQ7tgBrMOOjZq1+CbFAblXVzXCq
ItsYMs2TfYbX0LCO+xNudT57KVfbGZbiehrY2k3sq5Le9W+EC6V5B303tqbGesaEL5jQSYAthYdr
648Mv4V2qdtq9i9PJPzlzyt9OEc/0NfM4yjDGmQ41eFkiKrCGuIFIYCFFa+ev+ySl23V7EUdw81o
VoLKDOBPYDGsrhS9MHi/fsaec4aZTv4dOASBMBFziWrJzdoGrqmF6/VyZR1L8+0dE57CoiAICYSw
gIzJeY/qzEtjXhKPhNYXLLDE/vpeNgTqsJPSxPyFouHpxVx8ndUxy+2k1XyeSNjFAJxqrX3T31Qy
TPqiagKv+Gpac6QxNXAgvtUHOo+MhVDb/dT9yJwqk/n7wB6va0ZEbdjvunECb0FYvgHf4nEiNjGs
i93EPGV7FTSLp1P5D7AxG79XgrMmIoPz6b5uw72Tjw5Dhtd+RJsnWWJLvc7VtQmU5+9UJWwNiBtY
exxOUq/ZGPsONzzHeQB5D4s74SENddB5+EyNzSLgWCk+wQA2ZbCfxQbSI2wON+sdsXiFm9u1gUhn
lZRi8dHyzEJ7hKjZ7Hnpytml6YT3E+cNW1l3dhp4GHPgLUHT7cYK8Cauo1h7iFxvIxIGgppVn64e
bXHaocx7086OXcm/gcq6WmEHuCEdt4AIR8kInGBQmqyW9qAcMdiXyXyA3kf6iKGYexK8sNqeDpVX
tjhFJl3vLtnDqd6aUEw/HVsacEtz4mRBkfa5us5cADiR5nrMZKx7XbNaCkr84+LBhUmHDdP4xw2P
YUVNv6BMcCTPTUWNf7KZUQEoNvGbtaD9yD1AwL43IxLlo8lkyAhHWeBrXuALFAIecjzeKf7/+Nni
y9QEnHxZIuj69cGn7T45DXWgOGkPDgViJX8IrxO9hDrQBkFUvrsFYskoQ4IAQL6Amg7VSHl5Qhyq
OCaps6STw039z7bl/b9GSjFcG5Fs1uI8FwCJod9d5Q5Lz+L0CkzKKDn/9fkY7H6k4yjwO8TAV2in
ug/sleD7cKvx88eyCkpPLYDyA7m8N8sU0xpwisf1cg79CvupOBDBf0R1s9QSQH6SXABKzzE+Wr7y
vy5LbLfzexmdOGBMingg2XWWU+g2PdCqroikrfvHRyAeOK00T76IvEq8GgSivoBkHNELFIv04VYm
84lNNBsIhkhmkbfMi6fweXdht/70snebuRPvJQX4YUAjtxrJXfitB/DAeHMMb9ckeIAcfiqkceID
Fh/J3nT7vwxONndkQSxhppK0txcNAHwAu3wBS5Wwue3vi8AkXhk0tLyA9Whl03cTi0kpihZhcaQh
87z+Sr5nedLGG/WnfJ12TBIPbMw7I/TrW/m5cxdUt+0XdWH/xuBPWu23WGgE9Faijg+wya3iNhNA
U/1oBo2reQPsIqbYwIug/Zu4f0z24ClcvzEfaU7u9aVJroiT6fkRZ1AdX+ZyZ1HqIZyWCkjygfRh
5mY/zLWLuXFR6IQcEQx6KeetxYZQl7wHEXIWdrt6HSozlFLlsBKZvhpgIW/3Vi3RQUEOuNU9rgyg
j/+16whvJ+m5aZHAT0gZE+BAEd7NjGOt5RxE2EFKl24QfQBQZM/U8JZ5U2sMtDUILLAT+HG642Yk
xteXlS4rlSB5W0kH1t7RhaMX+zOHgNeMa4hbVV0r6LTnbXTXE5Q+JA1Rf5+V8Z8aIKSXX5Eli8TT
huqrWU5e3Qz9Ax8wWfmLInQEq6eOs0pIjtMBw58POw5xzDJf873pq6xHn+eEkkq2adfSAKR6PeXz
GhNviQ6UijIxNupX3sXct1Fh46RAIJKcs1STnouM1RVh9XPRbRsuEIXNx0dNE8+uNs0WMmyis3LX
kq9/wjNkaLIRwlX7u9dHx2UQSgtV33r9GSiy3yKX0qlSF+GEWlkvSDIPq3eSvg23825z4mXXkgez
eQfLXuQye7BMZ4MOLJqnbRLy37xlYzvbnEmfDbsw2XYXf70p21+zU7MJ8x1cr2fpRL+6I/JR8/Pe
WLeYZlFAWCKFbO4F3yNNMD9zfh86zEZqbBnvocO2DaL1mHy44yynlK2o09lOaCuE4x06Cu05t5vb
6y8wKqAg2zmAFWDZXE4owd5Rv2/9dFBCJhOLd/7FFhvCveJYNPRy0iLCKAU7bVHCQPweRL6cKP0W
MIj7Q/sq7LrKgnS4numIJh1jv6CWWrmIXct4kRIcun5APAVSIARSpwIvIgKn3I0vCJuUYyqebMb7
d3Kv+vDHgfd5zI9gwc7Ts9D7ByNovf7vHceyBXU+HaIVwW67TvKvsZDnFh3W/VLdvik0Hdk7Co+u
7ABI6SfxRyTjapJ3VnsWuVh5fgA5eZisFuiBnuwKzj03OGMP1sZtMbYRvPiyaVLjITJo6WkHpiPC
OjLkhNHX/HdUTifhr9/9LZ2nUj0+3Bzi6q6dQYzg5tE3+LAJeV2blNyUvG/wHvm3wjzuRiq2yEHk
R9efER0W54q/gkQ9QixIWbhS0pr4OUJYLpRGjNRWse8d3B2c469qXSEer8M+ecsA0OzbW81US/6K
ko5bnhPa1obq/mEIXPgtXbVzf5wdROZPzk+BAOk25iq4irRcn3Yozk/DD7yxJZwLq7cx2mub9qpb
S7PiUixY18fQgkTzvUQws/nIaSHel7wOLnN0ISsUcauFm1HXxQ3SND8jDPPJO25yRaYo3v4ssj0F
Ir7Q5WnVEzYqm319cYnxHh1NHkinlLH5SwfmoFqGWRlACuvJN6nDSRoDKAJd7L4EcpnroGvax/sn
eMKnTG/Nu1p7foiJVeMRItLS1lK78ByzWQOw8DwoiByKZ9ADDBnwVAvaPKy+62IBx3vXhjyKSwxl
I1jT20sznDUNjwCdFD4n5C6P7oQqIlFBbLs88PbTM8wUZ+Y4pIxe1Z2byfsAP6cgJcc+tymNExpM
+KYLlny/1T+Qfa9UF4YuIGAiqk8V/VyGtxT0wgSnJ14npl6qrzn66ZwC4cjzotJO/xQ8/L/coA/a
IH8v6BGP6sxqezL55aad8ArZtgKtVa1LeBoVa1P4RRYKxte/4Sg0EX286tX5k5/w0FVB1J8qAkkW
MulpHoj9AEm4v1dzdwqOZdskZmvppPVNwB31wHuBc/XhdHazvffjyUImrnfRzlWwd7d+sBYNebrN
UewW3TfUl0m1tY+4mT6LluapXgqjYcSO65REpWwsOUHFiPFpb1YImX32yH2QwW2rdiIoWsktQyW9
rbaJpuevIDBHdH9syeUxyebKScndTxz8e3RPYvEHl+rD5y10mq0EIrnlnF21/cAGdzgYgcrLNFvm
ctiWfQmlQbsas1xCuNfkJMjwAgV0IXt7QCkATFo+hb5VpgaSBDTB1G3iU+J8nIUCj/77ab2/Zvcm
W7da9V0vAlVmp3ZBNaPGu8exQc5V7nBw+T+vjgj0SXJkv3g5PRpp9iVw3wh2ItpvDvd3ZOnOqRSV
6mMZZiiHwzYSBB35A10QuiiEM/SqYS3lRKWEnisjK2UY9RgqrG/SGPXaSyqWl2D1rB/jPIkSI4HJ
CXtTpnyi98kvisljQ7nSPQEyOkj/zlXupJh8f9faJEQ/NMSAdSx5gwIAuYe/j4cTXq8XCjCrznAc
YS5uZdnvE6vUCwF/biNr1OZptypqRKfFtzl/aZOmh0ScPYjr8Hr15i9hU/+8ziNLZ4WHV5C8QLIY
KQLPivvIe155jsGycbyoURcC4FEPlislLpDdF/gysyO7uTHDgfLGKSKX8QQoK+m1ffRtNoPTCAIV
YpidSMEkk3+dlR3Lt57Wilv0RZxrM81yUDvP8kZXGDJE+QtLRKt7WQ4RJ/V2XnODyEQE2qsTmZFZ
HOx/As5Obd5Ijq+xuoqeO7OjMyL5kz6y2V6ImHSunuIZjKSbN1YzqrVZNjKV7ma+GngOcglOkGhg
Kq/OkoqmSZBFD7UCnwcxWY+sFRe31udn7uanbihC6rm3pPJJK2fulhQwOS6fobERflA6YQS1mzcr
Lqe1hCVTGRcYgP4B2Ej/K9IjIbX5zzKq8b2Z+wft+MfOco+uqiOs/4zPCMNPmx5QUF19swondb2B
sJRuqPQgRitlcOD2TjGpJpJlTawIaqWnBgA4DkpZSnEXxgk5jl/HGE6U19ly9McpQp7Ct2aZbnHW
O6qPHr04hEtl/n2I2CiBku2L18urXrypAp0k8yNgiNoEil5WuNTQ04fjTq+2GYM87HUFlBRYdbUC
wvETOwhILo+FGdic5jTocNXGnIYnYB9JTfrpFnjEHmxn8RXRINRLTO4JH8sxvHoFbg+7pfJCBrrz
uzCwr09zEeBWOK8qNo9lSSLzhVfz2wYe34BgOjrxv/yvqP8d6R2WsxWam7JHQnJhXNO9TcMUgXBU
gt2UITX0uWCvlOUEXGCaBooYABe4YIb1UV+jNPC9/fXjP5lvd4gG4r4BsJkiNpkuZxUiw9R7f75B
3e145eeev9HdSGXcjNYilZ9JLALlyQwn8c7bWwN7xlnTmfJeTlQHwPBybunu83oSen1TKt7wQRKc
hnF7AWBKp7m1hM5xUhfCRs9wf9JaWFa5AagjVZ+dEs3D5bMBfJ+8/8jfRc1q4MBJ4VMkXhmdvDIK
abIIg7yivtEt4cYpnkQLT4h9aA8kIxH6VRWyJiwQgBdTHhHt5d/E2QJSFh1+9qA7HhzWq6VjAmep
menk0D5pL2YISRHhSZg/JcNMOcjKTOFUFG+yVlE4Yl8/WEp1uD2/iAAnqKxQi3MVL7vRBFNGLTsf
jUYJrCtb/HJbqeUn+OT0IF7JDrezKFyOW0etz+hXQSQcmYQgVUlsZNHelQueArYaedqUeuInoL0o
uFFZGGXKqccNbnNvQCPbnyetX3HzyqrQJdWnEmLIKDyQEbV/Uh0jr5ra6jF18JlpsCcRCQFWuWbX
a7E8pXOb+lBrNGhAgLrc5n7gwbkX63AczIqmoj01vy5vshusvH66gtOlEDRv8YEolfDC3XhMhyiT
huxB++F+ltqlY1uD8jFsOTO0LbXdNLWy6cOhaoLr5rZzVOidrmPRGdwho0NGoqahdA6QsNcusEeO
MW+RMCWvxOWkIi3OY4UfsLmll7QdKKGR1wP7KiOCW6qK8XoRaTV6DFtCyoCpv7szuxpbsFmN4+cm
fMbRZrhgQ+jTOqOmUx0q8WnHgulJ7phXhswI1duBwPN6jogRvo4yzze35JwtYnCMzJkqXh9YIbx/
cpmUMZIlK95vf7jdfsPR15//WqKkIJgsOJEfR5IDq2C4OgC2SJBi69YBh0xOwL7CN3dgc0k2W5yF
/ZUQVdUKpN8gli4RNSTUhcH3eMHyUfOlglnxMdaP25hUlLWc3huOjkkni0jpJsKft8IKTikTwdfe
hY87c7y7IC0sdItiKqcl9HE/bSOwcdLqyvUVVQe6TCTkssd3H6MjplCxHxPaI9P5lfleCqN8Ne5t
YHk2ZwuqUA8m+K+Yg2Q8WMqSqaCmp4DSpQZ6GYM9pw6AedYrw6wz5HpjOwsmXFyhGQTO9GY/D4Hq
Cinx0loznYaUlXaTy/cmHPx4zYOWyf2zvDkvtt1fwB8sLJ7Dw44nJkBwQqj3/wKuSBeI7BISLKuD
INMNOQ7uJIuFAJLfvK6KcgAh8NgSNQIaCadnkdUPT0Fp0MhGkjHbuVcSzlmblsH0QwMRUazDFpvd
AIW1n1wAnoaESrIz36ruJczV6rsUG/DBS/udrJJYJSM1/zMS+MGqW+R6CSQAVQ4HifIg3uuB+eQn
HlEoRqtQxXnR0mce/teA3qwhCLDSPRmjfaXVgyy6DSqQtSNuwb2+N8yGJDnV6dZ2hr3AJJ5vEtGu
4zvPEECdoypEldsEOyliL0dVsw0vCUaxZmaG0Bdng32QU+vehBYhHyveYXQHMfmPcB6dtuUTfqJx
VITcZI9CIYbio/3kdjs0yY75+cCVFLXYxICvwTq9mhA8Fljc1srGEEBDDuYYfVJA5CoiaqJyIUGu
k425uawHkFlu16OXcClNFw6eFeITBD65PUUWMxQFSghgVuDz9zFSUu0waJLRlVJNN4QAG57RBdpP
hiTzPvDezOAaF78TWvMp/nMl18P4Qx2zWKHMEeUG8t47s84SsD1sjV1N7bSEBPPZwotBcxNvQ0Sl
ND5eCOr8bOAOnS+N3JnC6qNPmRrinQiI+a6VdhglUZCIbiKbsruYTIcNsogv/HqXN9/f0Q4YRZzb
QqWM8iKGzZRExQ2G3tj7MM2vAeOYPaUogyP58CpSXf8TBmryA1L3tUX1BOorrp0cvsfTbmG407O2
iJjyL7L/nYEWZ6bUTzGEwrYF9xtwmuL24SlDkKJMhw0JeA8Y+ebZuadRunJyOrmOEn/J8fn/4+3z
cbz3cCtlr4DJF0qC+QKrYLaULLJEsizI0ruMKmqP0F3YkWNUmPiV7MTPXQ4dvfVYCZG5YkpQ+K86
3oIrnG9Dw1Ma7zqFZ5FhL7Mgomsw8X/1ksIsLve4gYrb5oP2LTm2Yxm9bbmO81yFR+fjw06vxTCJ
hM9bsirkZRVHyVxnsAcNvhjehXgOF6FaCZQ0b/RDjnPsa9IPOqfBbB3C01ZwL3F696YdZj5dDc65
QNIb5PnL+QDazGp97Fmc/bY1KlQnTgOXsYKg0crRYoJBKrbXsZ0+YFcDj6oiQ53Rtblz7yaQ9MLK
8JYkle2taK1CbzVu22S0bgutj4EoL3uqETTX6pb5j1vEyCFSbl7SBS8XcQ5Hr1WrHQgwfnh+HJv8
7f8UnlI3UrWeuTZebErCxzHNopEzmWuMmkc7bDCvksxm9xqox/E0+TWjwt3N9394TG3VzaGAdP/1
YV0XACHAQ0phq9FBZ+SlTY0/Bt4sENFwPgC8i6T3X5j0SK6TLLVK3Bz+L7d5Vwez1zisY8TSpRcA
E+yhV9abMaXH2acHdDQ7it8dmyoCJzivTDCBjAqrK3Hnqq3nShG7LtMNyMUEnNusnbohev4NATuC
fcXOcd6MKABmQUePAxpjgFHZkCA4rwqBTbfSBzKa6ob61X6tp/OOU6DdXMay7TpfdtZTno3KqXP/
urnAkw1y9Kg/vDQEKmvhTB7b8n61lTDtfx9Qt6b7PzAmkhIAwwpQ4XYZOfSiKoJT1Eq7WAMTqWVP
jyll2iHAK7YKKIgtN49f6PF273YZjUkzjXnyJaJ0c2TRLuJwvPmAodyYzjQKtlxaPWypnzq7o0rM
uLsC8Xw4xbh20ar/JJy5gkIQaTEDKuNGC2j5AAmN6hpC0XBF6RpN2r2vftS6c3gAxBC6oGhJ8s6N
SXw1qRyqia45+wq8hllNqM/f84vt9WfChgAOPvaPiSmfZWj9VekgWH6D+YcXkp2GbNp8is+njBjk
MswYmeeaIOejwZJ79lDjIUkc7jHqOAUs1Nu7F/Pk92f+1fqKVVuyI22vgZ0heX/TEjmleT3gspGL
tpmk9QJuV0cg5SQE43gRppx+hzSkMH65VJFzcslgbdrAdt5RMI1nFOMe5lthiU+We6Do3n1zuzYR
62abWHgoCKIm/j2VBS6/RJB70pjTV5lZH9ze1um1o7RA71dlezT8rN7h0Dn8U2GS4u9t5iG4GOAI
7UUOHxqV3K7OI7/YGGQUzdkoIF3KoGc59nHsRNzoBcvSr4quQKXvPXThEiMdRgWEVz5flWqYMO0Q
H5BJ4CALQlRs2KGU4WlfVTygVo2/sUCb90D8sCFnK6HUQkepRATh0uFBzQ4ij1DpGQvNBO4079P8
NYUod9LNA1xnmT9/WQGiKDRo1ipIHk5mdtXA5VGQ1lGEFi7Hhz/H5Dnr+KCxMyJjO33SXx+l6kcS
ZMZxjq6V3YFVl31Tk6hrUxUTAg7O2rk4e4RMLumiZfdSp3cOHU+f5+kBeeCnhNU793cu2xgaINso
CMrGmMGcUSO3RQhSeJ6xJRDy41pv595iUsLlAzWbRT7Un2UZbV4964lwfdlnFANoZI1DK5sXEtul
JuuuBM3Okk498gsawlbR/gU+09ohvQbxdZrqSDHG2imRTv3wvpwochRlhiTvACqneDtdMOx0djYW
fGykw+3ci8uEEyXL+mOBz0QrVmEHfGIU7rvvQWpbis4mIexsvk2dDZmEzlHZ5zAmHaNgoSZA+GuV
Xi0TVDtcIzOGj2jdHxjvzk/xYDgi0cwGH8RRmuDMrRS7fqb9Lp9JjGtgv+50zuXUpRGk5wNY6u0N
YHrObGHw90q0eAU59x6/2crWxrU+i8nI7Uh1raeR+LJyNtM8MDOuYPtxdtbeRSgdpop2adH1v1YV
fa/cAhszJ+bS1tvKjz3GgIWnyeCl8jWW/J8gBQqboxWlo/exXDBbN1LWq59vv/ifPpsGUbD2VpFb
9vJxLX4NVoViFxM5Pxlpes2d5zSHrmbGY3VyO5fmg0s/j0K59Zf4MhPvdcWcIvVyEY7y2Fp8PXLN
potTSS0f8uujX31mMBaCuTz94Y1JLi3coCZQixetUrXbL6ExiAZ/3IWMzVTdJjMTAFJ/odhnBfLG
ccNppzhogVh3ScF0qGK3QcOv2r+TvymvxDv92R/0LrYnpHKnJxkI6+1iPudJ5YiDZyIj7tRxnjpk
I2VEN3mXMosJfhvjgLk86KtSpoNVoTZ2LGvB/Jj2L9xqoCrZ0nBx/gv3bqECWJI8k4uc0PVIQPIb
NCFEVqiZZzOEBM54g72UlF27A6zp08AdOz/GJR7TrE7mIcCB4pXMUMBb+WSDvxa+8D0CakuXnT59
MsNR2VfCjRBEb27+fLEilaX9QdQbuJkgVaRnjWHCj07wDjaWYDpzIfh9o0wslpfMXtTS1oMfZ8Rr
z2Uj42wCfdfbfkpLRLqf993pzeAnmZhaGcx0Fq1sIGOeDM5I9K1atw6l0crFEQGOUUzKwF+/5vrq
3opEz5aZOg5fKxlRg9AxMulQDNqx2ypVtn7UjvcKDc5YV195sKTxpgVuNBVqLPVddHb6wpjd7xZb
G0Xgq//7QBjSLQj2CdHKuFXdaGVg1oVXiJO5qFybebuYK/GtcukFIJP+0uTAUr65/pB2/ZXUKEpx
baA+DkYKULUO0YOv3gOrcc4LLcbWmI7qsLEB/EUqlSMmhDrs34xUXgB1aMAXUbL+P1sgBjW6FBj5
gKl8iD/tItPmJiA3npVww1zu89eIfEUmppZEaGNckZbGkXZzTrzBKpvkI555HY99sDOQvcBSzDSi
Zr7Sjb5bLHGhJfA3/3HNWb9fdL6KGGRedx3g4DD5k9/Yhd0rW45PEobr0hVRtO6prusdh+faMTIJ
KBdqvL6og0ujBzGcwJhU5T1iJhe2Yc4JIrPUuAlRwJ8e1OwfEl8VASgWmdGC+8ZOQx5GR3f6wEBz
PFacKqHT76a6AnR0M+opGtcl/Sa+aEgrxkJ4Kzrmwskems5MXESGvz1uiB05PZnNaV5i+4jYjMs7
epu7ifHTz7nRKGBprTS/DJw5QindMXyoRi9NjD0OzkY+paa3gCPhnnOObwOdBXPyGxf13AKYKFrq
7UnEWSw2fVFBeJoo65fZvY6nsVRdPOOhcamn7coHNDSCjFAuDYlHyuiJhHVfxJdD3t8eSqg1D3Tq
2x+y9j2Qh/2yxx8nHE0VAsNKsu8HGUvPYRwTpD4mDKmHTGEKEUmNMGSrh9ZwUTVxDYS0k7I8dylF
cWzRHDWPK3rEN+/y5Ls+b/74ROwWQQjCjekO8P60Vsnk90/sRR6evWH8PDyi4PNJuON5wuULRFs4
WMy6Lr59GwjY9S5twhpnAs+3EaO8bda4GSujAGg3guEneVtj88fsVMn0QxvC0JHwnKbdWyKRh7v4
5UGMUAAfu0PmbysVU2YktcJYS4VXi/5hUyf2k4ZlsbYphjasYYBYcdAKBCASSdFsX+FcpzMV2Qtc
B8+Fp7rfuWvaCwI1qPQmZSYhImM9j3sI3mvCsIkmsHwrDhV+0myPPUlGD3SRY+dqi2NWpnOlZIoD
vbWwJQi3Up9naY8XVKLNRJZsb5O7A3+bh3IDnVJ6akcYTB6J1KzdlpmigYlKKpkkSdChkJNY0ZJs
llrSwOLl+d7gFt6j8iJfumyk/4WpuVLpwmsxOlkhVFvRHvqPXnwdSDBleivTjlIHHlJkQXta8bvl
7/knKp8zbNU3sMOUgJXXcjiT+Da/qgQkVticNCXwZFwGC91ocgWrBULxEY4phAXKEclH9oExGmZV
nVb86OBGt+BcKA6HD2dC3KdHDrBf6XCfaMfKTGC6BJ2VdCB18x2Feqgz8AkxzWqp5LiXCs06dBTD
ftRe4R4xGSCiNB/yyqqmJ9s9ygxT1YcAKFUPbJMogOXdiTIcJCRKgg2G/BcK7U/NVC/goE99cyjy
CD0EEWShX43k52VDNw0S4KFRRxgLM+zV1m/XrPS4cAkiIY5KXHOVvcARAsM37eCljCLoJIm1qrou
AZMiFgjvv8P3PYB8Odk2XoWfJpfiIMcQ1slS0MqG7BAibIQRXu9IUBOOITVsj89T7SeqIwSioJur
4EL8U0ehBlKoj9GFMvfWgplMqadBsLdKLuL3800LurfRP27xYWLrdnl5plQUv4zf5KkKCmtYAKjU
Zr2jaj94HN1WG7vuKnI49evGOUY/UGGyebXzag7oJ/OPQdnyRoa+4/fIRzoNjLnZxLg1q5e9l2f8
4rLD4Xq71FeZHu/1ir4cgdU5Y54wZPiYzrWX0UQ9f6X5iCeFHmrF/6F6UOgu+ZD54aZHnXdoEfEs
SJ63Pj6m3rRWzNcSbZvu7T9LDqdF3K/GvgHW5KPdH5suojvTizY0iPtUQ9/zA8i5FHHwov0TkeCF
ugfwnTOig/O8s/3hPcaYK5idteHbXhXEHPU6+ZjX+ycYdTYBu6YBLKFMQ9+fta7C1u0EKgqX8WA/
j9EJijGo53VYLbI9H40Ap7lsgOcE+tZnHTMaIHXm91dPRk5PkUAbn3o/xC3IILhWr3yF1fiejcEq
QjubTBs3sPUCy+mCETlM8Dx1/HykxVfq3uSi3qbGpGay1N/H8fjTpF8WYUUBBbX7815QOdlPKigt
UJAb4oq5h4lxD9btHYutak+HGTcPfOnYNNTtaSK6vwfL+EJ8E/ZObQ6JbVY4sWzCXeLi9QfrBsIF
i1rYpg8k7cJkqoK3uQX+7WiVtfZg/hlJLZnUDqeS1ziYQqOCQTkGVuY6KRcffJ7wuh8ewle49lnM
fi3bu95s6sqbaPCEDoiTJ8P2OYGtHmbaexfdua/yuAR9Q1V3D0u1oOfUsODhPNzPSAffaKFKWGth
J8fc7YxJ0pJHFrdKeUj7j05lDOS1Lk7GV/QVsw/1FZIsR2zMVX7MTklGLI7CrhmD3Z48oY+kyWZA
NUUOOMnYEfRdEo/VLpuWsPR0NWcPuFUgD1oms5uWmr86DLoURp9Io1XEx14El2IPo9N4o9ll122Y
jiMy/Qcv/Sm5jX6I4fcUL1NzFimugMQWO2XDz48SjQS6mPv+Vz1lxCYe8H1RFZsXWuC2KZem9fsB
B8VdPDZYG3MBdz7V5jE5og4BpUsXIpA6LYh+sSdCms+jrCCtJ3X8WDy29vaqxMnQo40UXG3BrdaH
BodVZcYtrfdEBmR63fZRQk4EUem/WCyztHMIBpzFsf7FBisYldQOpN3TOMK04c6X6DVoCSOxFORJ
ZBaYnemBdp5buZmBDSfLRlRm/dyW9XzGSxrG+tmwpxTxPaJc6cbqcB37DJdv3qme719ElzIDeQau
FMHnDlHHwl8U/Hd3ZLr166R2FNs9xueSwzF7HNMRuzeHRUihLHXOahKeWzgPDQZlRQqzsaJjFZYv
zrvVppKC7pGytCfKHu0WmVsQaUbvy6SyCTlavYV3ZJVFwsqK8UgtcTjh0hXuYbrWd/UUgegJVsQq
JHzIT8dLLCHeccUakqv0zqLuXMrA8opRbMR9nYd0Juj7/EHsjhfTc/fa5oAHIeIbK/u+MXoWmBjS
Y6qJV5/dPrOBBoUJgFPt4trTXLotQ/cPuNfuyGYVzc/at2qi2al4xoNOIWXdaVncd8Upj+yBPrJb
UQZ6fQFOUOiRQXQ6pKIHDPtpupuygKw+vf99ErY+1y492FrOBAMkBD1KR1E1Ls8oVtAZ7ZyMHkbO
xLpHWyoQCaq8FkOSVYbtvMh4pVuujVeLOs6WuAOzAwRKDdcpKgMUnhpmK4mI3jOCpIi2C4Q4ERfP
q6EUp/piVYhnstHpkm+u5b99gFWsUTRswwnLlbLZR7bb9kpi2ra+raIpM41SD/H9Q4thiGzG0vwP
bqPxNd6G86hJIZ374lJsZ+OJvRkjhqU2z+hgpf/2ZRgOXd2KGhc5GbADP7zXc1GYH9VOkz+zq0LP
WNUrPEE5HDFBtVQhzofNkdm4SUI845se64Lue+p8lvCNBka03dFVV+bmUIpFM+DVX6ZFWj2yiUSu
rjYvIKvQMFNoyXWfgBRsmzdPHk2uTQJtWzgrc+Z/5KuBH4zsKdEXGIOwkh6o5k75oBvrs/71hpjz
J4dlJsi8FKFuEpN7oNglZ5L6SSV/qpIiaIXhPe+nb5QE1/bDcAP8FGfb5+OzzBt3L2zdVLnPkJ8s
R6boKgZkAdGxMj7+j+Hyptu37zjGG1jycXHsY3i6Sl86+wwWdX4iN/AvJWHVKX3wLRV3IWglIlW0
GiFNMnjDlHqeMiK6Eyl2be4GUJsQeNxUN4m+qSj2GRvtPBGFCF1JXLYfXVGkknkH7fDgc3fppTXs
KGJTbuwOhAkOFKyPh4HdHyO8sp1PkLiGxBegCzeuecoRSQhY11QyKDfHv+pFFEzL1h7M2l1wB96A
ht5Ro3tltlXZHVcpZJzfTt/efJbw8+MdLf39PUuGUO+DSnmhVIPSjRliJwQ7BqKiohROob1o8WdU
90sRyTmUylss5ufLG8XJ6qc4fiuU1R8x5Gk3C0tyOT/mLukd50rgy3UPCaU7unEFT8wVVOtb2+Tz
7bCnsSwyAc8Q1RiK7f0sHYujUK05RLXi3d1F22qsKXBDNjdJ+wq56b914vMRMcCO150a5kWGP17/
Lxc1Rk7Gt1JbVUU1fd8C7l6xoabtbP7ReEI3BO/NruQ5JnvUJjEXvslIOORThUm+pWchm87d5A+D
N69gafoMxtpQYa0O2qMJ1mPwMCkSWxd4JycjjL1x4N0dCnsQPHD7W0W/2cw9MewFxnVPLuVHunBU
79ABRIGZg8KjBfnp6LufDcHejRC5SSXdPQxGRr/mpFCRo1ysJrtOvuk68K8T1ixzYdBPyQuezXX9
R8zbGgcTIG8aoWfFdUHpmYypKCXel6yMLwD0iDbWT3BiJ+bK88FB4ADNB81ZZ2eviOzNFM2KppiE
A4rD0grLpiJvV7WqnQ47Hsxxor8N2oldz70zcIaUY+oUe3oqiiyExMMBJ0ThxaWKkbIvS5yQeTkj
HyqCJTHqbRmRQxa+h49yZH3w5Rf3oguy++I0ygBxwMPXJ3sVd3uptMCumDB2KiWf74HWmwlBh0H5
gqruKJEs+NWNDQCfbGIAZMNxdqsr6M+xFFHnWk0myJ282yaNc0ogelSImUNZBZ1o49upauOEssiy
LYUUuQSGTOP1nALGa2ivxI3dD4kKACXZg6U80CIzUKSMCIEGyohUxfoCtgxn2OwES/Z2KP9uW5S9
KcFrzElFh/IDNNX0AbxD1i3fxoK6MEEk010zbf72BZxyMV5jCnzkkL6gR5psvAGbNPyV2rwBAQis
DUx30h/u8hOtZ2C3Xr9N7aN3c2I+JtpGrDX91qLG/x7Hr751FfAoIxrIKS3Zatf/a7fQXrSy16US
SdA9G86q+IGvhaVd2Lh0p6jHh3MMcF/drWJr3G2LErJtWVH8wJWltnh7YeECMLcHIudfGP6gKRao
6ID6Qhlhl1TZGH0wX2g3lrPw8L68tJr95cf1SK3xtLil1/A5aXvFiZ0eHlMMk2BKmNqA37QUQEXw
0Q8GD4voLqXDKZxkLywO2PmZHhjfgiLIvZVx5aMIr+3nONv+gmbID6Thl+HjB0ggOWD9dlok+v+i
7nP+QFR9JazREOUt4IagEfkcwTTJujUqsUObJKLSsDi82IvSyzh5s9DuCPRbkSlhf5IWZuLh2sy8
1f32hpuJzrDojeYsBa3/1qpOHGFNw5hrF4frwuhQnTI/gesKLwZ4heJeY+a56nuprk2JUvXCzSqw
vYLgUH+DsmqRMg/sNddMZsoTxK0UpH0SVT6bDR4tuxGCmJrCPNNCsWiTktusxB/XKfzLp8VN0zB4
tv5yAIRcH0i/e5SR4enfJm3e9T/vp9Yuk6Ei77/sUhhyz6C1CLVDV5ZjOyKMdnazL03ukk/rAHwZ
JC0WRm4YXiV8aK+9/MIe3RUMpO2zv1yctCaKWGe8cgHSiHwjLKMS1Ozf/1teWvXA78bIPuAloaXR
utFJCfs+ny3sw20V48g6bukcu4VdK9xV63p9p9PNjr4ZCHR2V0H5Ih3PwW4gMHJR+9e0UkARSIRD
vyohLwBGFQhi9CPc3kxktmyvBqjDxQNorMittvIJ0vDmfzUuZkdnMuvNcPw9ArkcQbBblOIWT+qA
GFffI1ooawZA/UpI3hxiZQUek5AVvBclL15l3nSpyw3eeDEEiXqGcW0JIlN0iRANQ48SzDljxaWy
nRNJeyz1tiPSlov4ebJ22R62tbOpPVM39uu6or7MjmUUu9ZZqHQSB/3fXgsSkxkHItkm9+Vly6gD
OpuqxlKDiXfsWT0Vcg8PHK0676kDldwd0cqFDeZtHeTKvsWWe7281BIkHTqT31wgttZuBOy5Zxu1
cg6q34S0AV54D5iIdtR1UvCFMU/cl2NWvzCOo4e4okhYnIhI7IcV5azdnDlKleuoOILze+gt/sVu
vYwxYegHwHuwF4eS9pwmqyEd5U87dDZk+HZ9VvUOP7ne7hlxssfeZhUewYXgGXBVfYL+h3vtuqgx
qaZ5VGymrxX63iwqW+hAjI+a6SFNK41C2eo+fQQroyA0v4LMTme+rm01zVMdBBHGcXKUi6eb+psy
CDOlCQhaKbSNSoIRGGi5nybFgsvjgNk5HTfUljZq7sIo/JYJ8wfyOY/r22RE+GAsSwJA/fH6QvmR
Y9PWnL4jRR1eQOsGypY+mG51ID8gUibxm9/kQG3rFuCEbBV5CwK0os4DfBRPkObssglb03EYsSnh
TATmBSkEdmBh39O3hu1xmlSTu5hZYqS69y4lFEk4VBs85mD1dJaE9a3IgJUCQvCSNwraaePGnrCF
PisHl6bwnQ1WfTArKdqBch9MXN8MjPb8DxiZfS5u+grNwxN+yIPTW+iEfyTCi/DiBuQoxTLjkQJ9
4OFCLKy+oXhYJdZdb4burlSMsFTTTuo7fk7HEM0R8tW4uFqyVKXSkIiQQJfgUO0sPyuMdrAnHSHo
fM3XPpM120hysE4IMfCuAlaSIZtlwDcAByq3FuLP/PmTrAdBgr6uMOSIWgmmgCw235Zp1VRrtTQ0
E6rasTxfa+8/TwJ7bY+p+MNwKptkaVsPAXt+yXzmSwQXQ0ZWWvL4hJQSA0dgpEEtPX1cq003Smzj
YlDAXiXCDER2/YXvFIlWrVRtZdFABFKv9zNUAPHQU76ytcFyQfhkhezsFbMFRhz0y18jFVj/AGBy
7V9anbM4KOB3Hv5ujca7RyN6cr7Pr8oWk3m/cMkXEb0GkkhMhlybIJcwCky6S5WUEr5ZvnLXTiiy
LH6eu+2Ys4SfCa8CclK1S5sqFq/4QwyUv55BZVTdFC89LgQ1gfXyTwrB5Vv7YIt9t0GiKoviYjAc
m/XYh4XuXfCi3avvLcb2+h2ga/Xsr3v/n99Vrmid/hVvvI0ImVmM0jk5pjW9kzLz55WyNXHsVIcH
qPpStWXgIasFTJFkAY6sAV5OIgxy8TAIdMiK86L40aOoCnXgXD1oH8u10zBRCKR3STsH2tIcdW65
VL+aGmu6RlCiSeO4pK2q5hs+GxXDAtLgN2CddjC0nDGfI2hwmqY8L3NoM5PVsQQUoW8W9Auic35y
5fbEbtMezxwnfiUJ8gjsgS4QP8+qmYXru387quc3LGMrAiYpYO4P0lWu5Z6iGQ1ff6Yhm8yr76uJ
babgP8T20J+qmJgaLCcYH2SUEwAVS9le6rCJGjV5qzSUjqNPdTcuF8xAJmy/9koz2hjRWVDz0bEZ
56UqxkmaQEoPRjR35Rk1nVpjBROJJ86knaWfcJwXlPZJLG0nM/kX7Bdc4KTlILT6sQP0WsFoD7kX
NFh9VsbnXOogA+Y6PUgUbtpb28RGTkVM81h7IENqlv7hzpHowdPxPMNW7Y89p84jySkLOIVYedpR
GFaWHfW+MWyxlbkuzzYY2pG3H52/xMjaK6RT5MN4ZMpgLI8ErpK3WBodURmdnAJVrjmvr1wLAkF6
t880Xu3Z5B7MOwZVFK+ret85cUCWc61X5QfG8u8re8ARL1GhZlzslfGjIF7jGjBjP/QuPdCaizvR
igUnT+h6b7NRqjB/4MRKSVXbRpprdnotNkw4avuYt4n9BzCw+OW4lcP3+bbSJnBy4UiBw58olQl+
s9ZIIasb2pBBJHWEHkEFNl1T8GbJqzVDlfrw3A0l3GkPV7Ia78IIbtkKock7l7xRjWt5iCeyewWv
EpJbCpCPzuDPyczU2P1PA5PL5MZpsS/4DWktZkqjCivv0buUNJetFGcCEVF8QJ8KTorEPk1g6dCV
haqUZvmL2QJ21XjGt6t6Bs70SaUrU1ta4lJ3hblrQFTxac4tcXPpb6A+g83u2732pzJEZuDBJ9GI
IXlIUaFT1VDvkBy/xUKRabEHm2oxy9D1x7jhDGwl+HcutJtOCTrUVS79nmJ2+ZsKtoHFARAYFue0
aDTdGCnoxKhCtwAYls8cMiTYDrcOXH6LeIzGXlOlkwFUsaDoJ+8Fk2hPdHCW3e6uX0tC3WexioYO
XZCmOvi0xirzqFNVXHIqDoERPzsu/6mOgEbajqtbShD/1Iy60Xzv4eQSz0LvoxXw3hcfO/QzxtO1
WRcUhEuw55x9+wjqohcPpfVSYIsEH49cBMCKYYlb6Bzwo9LAYVaHjJMDQQBbLPGb9Y5UuKweasPC
G2crY4H33lZPTbI/RpHKAkBTd0BPJALS6zNGjiMC3uEggCfQIMjgpsc4fm4wo4X2qVPtaAPYcQEm
RAOAFoO7T0jWzXkRusu/LyLfLGtXNXUn7XV3tqI2/02JnBvqqMoGO4ZsNrhf5HTLYx8xKbyNEtId
ZsMFQECNsft8S88+qnJnKOhWDRisWnLg6Cd2ieIAetsIeX8b5pDoCoThvScV+BfLeyMURUCbT6+2
pTAsmYzH9I0m7frjXPHFqKz7o1gmzgXV6kJNMlpdwrMoxs1TmeAnEjrmt1FuZ0J+FeDE7jwRNa/+
6lQNEeJ0b+2Wnqe9QpqLZjBOvjSEqbzxARV9O5vQ998BMD0urg1nJbc3OY7hDW8GvUOoreOJ3S1q
1UFimWEFeDjjw1Latd0m59wCC5mDmf0dqes+ccQs2jaOhsItO5DHofqo7TKps/bgUQzk4/KfKElU
RLGLua5SK1eKrewD6X+UP1FFM/AexYLg7+2+gbNjbc/p1VmItrdbVrMQm7AugRSWnV+QYahLr0eR
gbOXmw1C6gijXKIB6OJcGGL7BG5cq0y0ws3il5g5UUA2zLuRAYrCj/pF/ODcni+LGRbNIDR1uYaB
WHMR81pa7OQqtrSvgpxFc1Ev3mvnYUnNs0sLVj1m2kzI/7ZvZEY6nhUU8rQfhIEaySh6V5lkCUg0
N9UomI1tq1vTIbo2C0WakCvqrnnbG4DV8ZoDSHqocYTdccvf/GixTQ/Di/8CU0qLcsvNUbdH7LxP
ytACG+kDf6EHPw83TdQfazSvD75CcA9z8V8aiq37cqTmWm58Nis1zHudNGhdV4GVwWwUJYDAWddT
6tbzVhKc3hs6ywb1dmMzojrKFncBYZ4h5SpI1ihGSvlR8/Ak5oF2zXPpp6ZgjhAWI55bFqudbqVY
DxcW82JQdcXCUfiHHxbBKEQ57DEWcWxMcJ+5ipSg8Ynli8wztM4XOpzYrGVPwUQA3Wgp3MUTMRnV
P+jkVvwvHWX1qsLh5hNrL9ZhI9n9CEvWJgkcKz9DGYzMHzdzBmoQQNi4kGCGcESujr7MKanKStwd
PWs8H75+Pc9ewpT8CGQwrru9CWvzi9D5/b9d/c3ZHVaSSQu3B5tQ+6sUzE2A0qXp4moUjpXkpSxp
EsMGRXZm+ZLBbTOLIHmpNY3SPIu06Xan0mlXK1jon6zJhC/5niearjTZZQ2ik0WZBKiK2FV9OCjw
7KoTMUxYhMHmp1WQg4M62Jd+3+WJcOs9+4ELuaNb6YJ6bqr1AQM9307gL/UTt7DNs0UbN1SuQT7w
we9Y9coFR8lnNUitxKL5J87PSyrwCGE9jycyogSZw1+9+iJek1Q5PgxJCZTHyye6mTl4mEQW4otB
ZuRIjIVk2dxgMVzqMbz3nM9nF3DBWaLcd6PdneX+LTDZSPElNb7nvGM7WY5lwE+bDHFZ6xs5lSj0
iOIURwtSNchv7Tsmu9pFSogKTPHN6UaPJYDQoyDY7w1ZVIZ3wGmZMWoY28+TzzmQD/YgIyqd+EoF
E6rjyhZxgRuHETEZcURKamM54aPo3TstWvaVumgi+JOkR7XrBVKCralpk9NaE5lnS7eY5tg6INhc
uC2cHmHFIWvlECGfOiz0XuSiWIvSicn0tdeqOgjUm9yDES9QNyi0PTMVfE/oH8eA7tv92Gl7/MnB
/ay86sjIKw2VRN5Dh2vfiCkV0mYzBqDOy2U9223W8C2DOZXm5CDPZoDXq4/MaTMxAVitg9//opJ8
vfXa1dLBMXOnAwjJotJgO+SpdyA69O+EEFfCezHOkKK642SdzSsBrtQm6f7aBbMwYOjokPFfnT6i
+yhbaomKg6R3gzwyPb27H5blKSkGC1byn2TSIp2UmYbQElgt2LvXmZ1P0sXk5H9aii9K7gZyrTnJ
VoXXiMTiLjMoIUEnM8fIGdsvoFs1sXUvyvWRDJBLJisfLi3jBb6RxlGdmhW/1CX/cG8IhMrHi7vu
YofhZMJGje82Kp4DzN7PJKZb/osHucTsy/S4fqj5cIkKnI+9RCv2EY0LcZT2+Pqvx5c/NzSldGL6
BzKlayHP61IxCvzCjjNxG9BxRU/KjVaKp6MeLfm/Zg6acduV51ftT0r+WWLMuN+vkiZh+hhlLWq/
cJAGtwVQg8+4ROq7sHgi0iISBfaTMpta6rFK0bGlv4k0vjpPbExd0Cq+Vr+lJAODTGS9Cawe5n4w
zjnppUdwKOizdo0lfFn6OP8pbya932bHoJ9Bc//Bq7qRD6ayN9/zr7iXTLlKtq9BFsDb3+qICMx/
3GlEwI/vNhSg1QY10gRlsaC3ekXyxKgGujpOfVLbRYuN+tZP1fKC2svSTpxDwhbylswOs7HO3Uwa
q8ns4BUUF1IMVBgG53E1WcK+pc3NfNhBqQWTkA+fiF9mynnHqdyr8+lDsffy7rxQNY0w1sUSIFet
8fw4PBzJMr481bBvQY3aFL2ch72exwjzOO6ND3qC1OTMzYhLZJIiNq3DoS0Wf8tT1iQmPJL+wj49
d+yQQiiwL7/b3dm+jZfzEEXGMJQkko3ZpmSqLLBplMSdfTIs0E+IvXs/tKTCv36DrXipoL+nWt6C
kdb0+ihv2ucTdwndzo5SK2cRi+cMLmOgRssMjaCpTSKvOo6V01uluvGPSR7zwo2pQ5RAm6hHrywt
GAnhgklcEalHDwivzARqVSVBWKVxrPpiiUMEVrHbsBBgyhP7eCed1RIDkT53EFx6jihthcUnRSwO
rLP88bIuzD1l4pPDGpV+mvqyW0nD6sNROFQoYKGUmNeGSUiVV7Jlm+vgaMWrQDkyAKsOugmh0sG4
U+5K+TwxLrIGfySNdC9A3JK07RN2bKveEEiYZqDcOw0ZDJuGvtlI3P+SKkKfUP16CRE29ApNbiTw
NswCkuR6/k/OSEH1JDdHUPCwu87oG7IunotplTqGC7++AY9AKlSBRavV2x0w46XVukmS1YeBVeyQ
J7MxMLtaxpu6ryZMYHs9PU3E2SJZk6XknkCwXkbF4Tst6ZCXuGaP/aYihJvz8QMnKsKDgzxpDKd0
DsWfc18U484Q6Jw2u0sPnXTK4g4uTe+2uprbl5W1uYt3r2YWXBn2ElnG05wjrchJZSYRZgH5f1H4
f1M1/TqGJaMv7GJ5Dj3dcEopNJbRf7hT342PH1JovqB+agAhMRddBKPD8afrCjzYFdNlp0PAKNrl
3mYFrZV+Cpzyp2+7eZSwXlr4MSIVBENo/CyX3XcYvRif2cfyPilzRpG4nGzHgY9KncQsQr/TKqQu
4Mt+16uWLNV9iSKULSGsZlAUD132Duw3DXUigwGQgPoZuAqbrCOtky6g9GGuAfBADB4IMidkmVa+
LTg6U9VNknfvhRuJGvviBKY4PdIa9Xbhd49d/o3CQBzNhgfwWz/H+PcMLEo+HDT66O4y8SOZ29im
kJivCOI05kOJy5C5Ppf7K4w0qN7ciu9GyErquz337SemvaYCne+LJtuGsH3Y9lk1NqykwFZUycUK
VmfpxJ+0n991rxpdZX3cWAhncvCSxBi1wNQRWJarHQsP4qq5JPG48wpyNy5tu3+w+otAOMkvzT3Q
XcKCXo2lM07+eYuXqQFfAP1wUXsjQqnafo2hXkDlqz6Ol4UztuBx9eqqIXK7hjYzIyS0CquD5XB3
2eO1c5JIbetVeu6ZsevU4P1pBuyahMnY2m0mL53ouza+xCSwVaQSXMmKqa37crdqkRIJRkBzFfXG
YHGh0gq4sEPnksFBL5GjjMfDk5cpdByX1kIXNvhuxqbPGfkGrj4HcwimPsUj0zemzGpnc1wL90hk
6hZCTNGE/mMhqypMhdWdAuv9JWaiUxI6J08v9rBdhpAjUAE/30L6biSDIq8rQBMbI334RAh60q4U
xeVHAZPaJ8Eq4eN1Hfm2VioP0o2GAKMYwZ7VQlzCHPOGb3ytXL3wo7aF+C191xy/fIREFt/wWzM4
kvlqL5XQGbg51xa1LBlmAxt1ZR6nrWIx0IyodxQxaD8Rx4+zTKV41hoAG5paJApc0LO7COZVWTe8
ObRR6+vmsS4s3GpucaFMMq2xf7B9iXLQs7lCbN8x/vHLcqIn44nZwfcP2Hc6XLCdLHOiv2tewWf9
n/Xw+Esi1Hqw+cEYsBYcFF+bNNRutGTlrZ48LJY1wK6wPJ6k1xpOh1N7+k4NRVGx/bp5w8IVKADe
4M0Ow/PC5XsOMbj6ztT69kM+F5eEs7bew3DcFPJ8uP2Z3nWgQLBSRCeywfORKrsRG7DlQhQl4LN8
3UogUg1HkNL3s4n28CRsPMborcRiXfV5ip/WudyBESpleXdstqreJpYcIXfhGa//vCvCH7ubN4jX
9/oqWe2xeDXd9IgVoLwqOq9AafYWWhn+OfuavUzUSfIDqubVMGTq8mb6IqigQ40B0vxnde66g4j2
JZMeMFRoWDjvHcVDkp+40ANMDu4LH/sWVzMWdYLlWOpky4PsoRrOlrtTxC4XnJuyAsVZ8Hmwu+We
iHoU9rKrFwCNuKm9m24T5aAiTmpKi7ipXNszgs4bXppJoIZTdJMX/lEJGY5wNRZjjDxTa6VjZXM8
rQaEw5phkatNmcvfptXPBfmZRddw2n3mXLKXYXC7h8/pt70EgqRmEHD6EbHqU7Uno8qEOToWVPuz
4cvFqm9mtvpzeRyf1veh7Ct8JKPSBJ05HsSB/GcDoTJFIE5C7VPqHlW56gXIVdrlJh/2GGNIkkuN
Y6kP3FT48JOgT1k/lmLWvQ0878cfERn+3RqFmHfFMg76juXjNkB2IdTwDxqCxB2vATaCtXhQiuu+
ro/YcMe6KoNmqHvERjzsPfYZBs+TQc7cFmoLvWS6PaIZhCu1HIo0R2jgHpFI7rYa1OxPr0avnwqB
ckM9lFPwl4xbu2dVDGh8mjzsNMdQKW91WF4gbPv71cuuGnuw5aEsju3AuMU7qQqYH1ZoLYwzQz+r
bK7ZQ8443uyYRIOdq65OLn8a5/oEv0z+8Cnegs4jFp+ZlkP1hS0lC5vdG/6admeh1d3jZqOkqsDZ
0ezCYCAhyhOc+AD8uFW8JYN58sLpPKio6csqfAFXRaB1JkcocWESgf6vHhUU1O1a7ty31ztdvK6n
LuqUKtuNkoSar4gE/BdxyvKz8y9ssKroyNUmk+fSRJRkSNy0iRKakZaVYujNiucDVybO7PXV7cJA
WBZohLQgWGEXB+eAg47lBX3Qrf3ipX5SQmpjspIVRuC1dKHwTnfPDZFzrntgSKw2r5ZGUjIBP8DD
yl3/iVWKSE969tmcVMur4LCR3o2MhklXYBlIzwcGqDvxC5vVg9wTK0l28BNLyWumKkAWCkxvJzfz
plfPWWcSfBBHnDD8WnYYHE8soN1kgtScpIaeW+h4ldFSR+tHTOHLfXi7+fbi5jNPL44G5MQNOInt
SGehZL3q5VYdP0GWx+MyvivETMoo6Ro8lpSNH0N0BlYC8a9DXdksyJFRQSe3EW8LtUwg1SeG6evn
bvhtmtg8DcoL12BIEXsZ4XzU4S8ctIghSDa3jdSL41Gawu3BErQofuyKMigrRok08RzkEu82wOP7
Xi7r71NhCrzDXL9pZRA1e/L5N3aX3F9ndvuNMvt5m62O2ytnxYBzI06lKbK5amG54D5KQgP6nRut
uO3uz99UpdpWfaNEk4EBJpzvmw9iJ73hwJ7Qoio6MrEibaRNYy50RTp4YHC1pmQ6qDwcP7unG1g7
7Iz4vqVmTiqnPUW5eDYCWFYVqjhi3SzmUjpmwk+x5TofFnra2VHh0nkOvqcZp4LErum/UJ1vGCyS
liEApt1DMT+ALJyKaQ5ha3EW+Y8cawh820th0aLIguGudSR8+264MszZiFOM2VKxzv8Ged61ldTr
5sU6klaqfYiwq4AyN0MetMH8RMMMbS4FTZ+QW43YSQVj+HODjaAe4ugWMZCiF0VDiqO4Wg0wWKqZ
t+WyaKaH+qsYm5qdXNTEXbu2PrW0nJJge5MsgLn2xoibO5X9w9L91kV9ZZ5IH30wREls3MIRYY1O
AmZw/VVxcesir8RzFnz3WKI0VSe5pXCZ6/1Y3kT6Xnqp72mMbe0mt49TkYqUEsDaq45by0xWLPP+
LLA0dgghXGjgA55EOoZjv6LfSpF9p4s0xNjhWz8R3+5oiQVbXpAMsSAQfuS0htZxRSYa5RPr0d4t
FNUeQahe2m3BG2Aaqo9EvNS9PgE2a3bslvOJZ9gcOPjq/cGNQXe//LJRwxC+SNTLAfafjbeiPfYW
OzVKeaDeO6RW9VNEqKFv9OLWHsDSptKVFnuYzf8NsecTxsT6Wi7QrbR0Xs/cuiqyMz/GcNfWtzcl
dFRENPoLOMlI3sLiRcvzCF99IR4RsZWojiMCVqI9G1DIv+NhsEINdwx+L1S+SGqVCmDz6F27A/VR
CRKmZBpD4GNjH9KWt2ROk9d0KEWHDCFpzNJMGt9nlVd539EHcFzHThxsf6rrWn/fs98qazzha4DS
iPd8gZbLbFzqi7iA4BC5Io61ttt8qYk5QEn8J0JPERNML3C8ar9rEwRvX8cegXQB8PLLIqJ6Zjsg
RHqXlPxETF/Hhcnf59fJMIzJU5BJHk03XnOjsszwFx0XrI41Rg+Bn7XRIhvkoS47x3DOrJnB7/Q0
j9PB1Y1Pknmj/bGdEZelLDU0nZKelnrCbHKjakcWcZcJ61DFlqjApaZbdW+KZUZw/8vuuZ8IdN9L
5FPnYFmY4Jr6wPYCoNyx4LiYdSzuZPYIQddsumBT1HWVGhnQQpr4CIpe2aNpHJcAKWRQAHIjexuS
+nH0gkmKVotGVY2C1A3YtxEiFMKnq877c0JxnfdiotIL1LyfIQUdcS098VhFoCOgBJSrL94IA2hW
mBN/rQ9JBbwijLmcMaud00EcitoU4AuJACYJpUhavGsADGO6i67cgRJ2WjzaUuZV/uXAEMe2QxU1
YEQSdR21MW53dnf+gyYbPf0LbulDVUQsxbtQJbqYgKj3zk4N4OlSezJbdfaVdrSbdBPh3W9LRInt
2f3dblThV7ZsIjHB1h6G9gu1/BXyt3fZPHH+H/EhZLseNGEZfvD4usO4Q9e+sdqcnXDA8kRmz1u3
XlRo7YsKhcZByw2eeDgZHbESs2V7E8XqBtAamUuOmkG3XRhBo6R/kN9Ypo8HOY1Jw1fqPjcUOSn6
77W0kqyH/vjGx/YNqoO3pQlEszh2zXl9oF7t/uLU/08gwTVkv7UOcbMgUdRboHFoe+aaP9ffm+kK
oZW4n+z6Jrt8g/gf44j+Swx4KO/PfWSAzVnZ1YRb4LBj/5Gzwr1iLOGVPmaFLqpZwUoFywUrzu5q
4rOl3ZsyxX9LS0PGT0Za+WZccRWwGwDfMheTWUQkiEhNv0DeJWnLRsYtLBTHxpYIMHHGVgdtgXiH
z8rNrMvRyQla6b553WX0380eTD1k2nVC0bXHh7j3BMJuh6NYiJvN2+qblerllZc5WARoVCEQLFZF
pNsbHvrb5eo06b1aDhy4sWfNRRSzKViSVIyZkHH3rmtv6HmFHRSbw3JNdAWRgBBduA97j8kMxKIb
M8z4cfuc9oxN2SV029p48HroScXO0YWohZ1ALLGeOXaS2j/tzoXH62xUfx1yCrCX8rGwsj8oFXdp
089WJMXz7YnmAQXPgEbjeZxm9e0PL/qjbucYVyd0LzReWI0IKsIZEADBxHjn5+ATexKXwxXtoE6B
Nwu6VwdhBL5J6TcB8whsquNehhajZIKXoYMk7oSQXQLi4kgv7JSRGmMT5Fo7016OtQcOH9Akr9O+
xl6ojua02nUmozb1XXgs3xPBqWxEkSCKPG5T4WmkMnVjsXDOMFtUgNLqhgnTCi4YFdYKPnvb74/2
aVN8GF5WvHSyD61HG2CplwYsQSE6wcR89TeHynAc812+tk2/SHnuqEwREA9JGh/wbbh9K5ud1uSj
oLVj+2od0aFbHze7dJKNu3Rrcl5LQ6IDWrarxrBhaTIff0dP4J/1JKi7SNeqSics+3kkTMy9vJ88
HIL6MIpwd/1WYlyYLRLuktlqTjzfMWfCKJVYgv3weAeyxalOpBNTWbTlG5AJTMwC0AWnS1ZOcnO8
pWKlLFmv29e4LrpuwldyR/K120/Ba2Njmet33iV0Rt4Z511oqNgbXs4m2LMhMy2yw2cBAAnnG6NY
JFhRd10DftFKuzhXiOTN+cjl/BANpgx/Rn+RjYBkQFKsPq0GTww3vQ5O64YpxzJLjy3PTlZXFVRs
7mog9UWaRuDnkvNbvEwch0YQUPV147D1FE+qS5QisTfeDM98hRnzM8XvKqxchBXj6ve85ATjBG/4
bIF7tryFkghKey7pZJ8NQBXxc+MVWMMhutMqjgrAHr6/Rx7ON95LEfVIPAYaJXQ4M4tt2PfdDa8l
fRD4Ca3MgHnypUSIKUpFeUUqvZXs5h9j57zwmtP+YowJl2Zod644G7FBMCRny06OhyYBAbXnZxf3
LSJL51YePCCtlRT6U3NHeO9PEn8I3NwNcWwwkX9KvvlDYAg7Cx0vcZV0DzDftVFMu7DsBMC4JClz
l6zPebeDI/Wx/kKIaEdNIrh0dOIpciurvwXYCtfU6VSq3pI0qubooLnv/B8j+Mu8ERKNXbUj/nkD
IgyJ7J+RrHSyQcFHr+cgoXycfnCeBG3TMnhAMl2IdPLm3ifxfsUohJ+dhLOkleXl7Jx2v2JSGRDD
tz68s5DR7/zgHalZFQanrpH2r7z3tzE0DjxkKsF9xMYBF7neR3Q+ZMmfb0/2wc1rqdJU8Jl3uM7U
+yy0mIiB7lH1GbfJh1IzCQ5S0TuvjOyD+DHP0W38PgcsgBU+dGNhB0RZ3MaEJbK0ezB6tmS9LT9D
ubloxSUnfn0zkZPJTO+MeHMFfkEgy0DnhrYT6Jsv17PyP53TOMLh/Qw2wW73rCPtr3GOh1ippUEG
myRZjgn0CuqOpYocr3dT1TF7LA5jHTcTofdlUMKEaOMiMkuATZDJ41nJrnQLTn8mgRDYt/zl4/iw
AX9Ojuw5y3OhnUGgXHbw6mJwVHNbr9sIA5sSV6bgyTG2mP6xSI3rJGgf4T57qWSlUBMMAsIp6ZGy
UyKBL0kbHLDfl5DF+gETJJKW2FC9VlQ9/DgwE/z3WsjcsCRFJEZx/cvvxpsoQQgWuYZ0/DYLK+VD
B9MjQPAv9Kgah8bD31siP7k6Gv5Pr27B2dViXU+GqLgreusE+0bhxWqH4Kt/wO9Ut+QkdLveQhve
/T2EV9U234EH+xZTjTXTBtvXJxhLndaCl+ejy8i1yUubvGNAnNG7DdUJ0cNdTK6CmbTQ5n8PwwoV
0tlyTkd+QT5xjjEiYI02jZ8C4Z57ExL3q4s381kmfveXol2aW5O43qs0vOpe0gR71475EmUfvax+
9WzQXesYx0fIeb0EI5XpRHY8Jnr/QIQUQGKy9BM5wIS5ni9e+I/pjQtPhU9YbfSJIYM7yLhzhd4n
e0zCxyZhTPEf+08gE/0o0hAeJXp0C8VBl0Xz0mEirQttP2Wbgoj6WLykiYXlhG7+/I6Ur8dePMsl
Z5zkZ/y1PanprCDDqpHIsD2QjOsUPzkNtAIt9ojiko8DtsUGLYnFNRFsLgyr/N8OJq/dd2y1sIn4
JQB+XgFMjvM207gnZuY5DR10nF8UYvrCXtb38fDKAGgp6q364eE2qJ7t5Ga2za+vqCWu6yFbv4RF
ErhMwjPYlGXUIr1OIFtG6eQqNw7LGUOepBoGDEQsNCmzRnZ3jeiNwCjcUDBgE5yZ4UTKUI1u7Q50
Pc7Zlhw7rxexGmYQzP/daVzVxitbuJNYuWGk/zxqUJ6OKYeF6oBab1zkpYR3es2Tn9sDbs6DAORH
5gNrI4h6Wa13OCiYP+PyFcmBiFPPhTqnOswwCGE4h8LQQ3UE1wnrqFqnrjqfsmQVxXpKiLSYxx4n
YZIVb2s6XQS00dce7fdzxGr3LQDYgulVlhqYZ3OM1QQ/yOC/YDViDks9PLt0TuAvOlIZzUR9uEfT
X6IspiLRN34ej8s4x0yho68p1ZhSjMdA39n9dZR7Jkr1G0ltWQjhaAwr8S4nSlke/VLaXEDlMp/k
moGR/Hn72ZxeW3JCNH1qu2mQ9o2tBgv6VHI+QX4BkP4fx6GELhqNbYcRFBdxdWEqI6/+2s++PUZ0
cyxZsnIVg0BU8qdzFkON2l1Bmp7NrFwkFU6JCUrwNCLjx/EasCJ8j8Y+yrlIc7s/RwJO2cgktA3D
bGCrovvfA9dxky9e6jEcNpZ5qJIjrzjyZ2imAnFxKe26yIT977hiOJMOd4muOTBfUYI00YD6R6MH
ABm0dKkEgXH5aOxsyx8wGQO6Qjt9R/INh8DvBiGhGt4mm0zHzgUfsdBTrNLCOnzgQJoo66n44FOq
PensrUwZl0CPJ0s+vexGDy1hg+EppQQTtrul7nf5ur+jPByyASpTopiEzoxrCf/K75DemYcaePua
zkmBkIB4vt03koy9K4VJlUmF+S+TJ30/AkN+kXeUfQSBy3WVgHH9631k0ChqJB/9pZj7GfsUDtJY
TBKz4Mwjn9zZM21CtOyoADUxU5mCz2UzsKT7cviXzawPYYckuQrNHQO92IlX8TiHmxR8TCNhiiTU
o/vvcY5XbcUDPoopx28jXj/V7WjiIaOT6+Vo+RephYYBu0fUX9kFIEKEKg8R1vf+jgV/QhNRzRQ7
C/pDP1i37fcYB0+u1FY39JKDg2fTvMudTFjRS4izkqC9umj+TkXUsurtyp4/GCzjgi0+fbNw/phC
zyt3nfpfIP0iCjNkaSiOQhhh6tWBeYAn3u2v2asoHVr0MuEHNs3WFdBggKP4e/gFfhW3GdAiexwn
OTuttohWaHosHPBt6VjPPu1xr8KVW5iXAlQpvqKNTJCtnzdFtgFkyRQszKijw8expoKWhrei3HEt
gL3me0h0MPxey1PJK8W77tVnwfzKJ8FuXnFSzVyHFbzGbsnWIwzkAGKE5rzeNFTRIhWbBpsgJhZ5
U3aH265llFwMgWN+BfsiiS7Hm8VhYKd39k/P+fQlxTeYrDOWTEe+KydApkY4gv8TfIzHE9UJsE84
MrKamYDhNd4s1cklThkAU2aiENuIgQxQSs4EDDCvSistipWvOshEsSyc2cmOlKcHtHdIMlfrGRL9
LZ/7P3L1LPo9nOK89AlVJD2rF/PYNhXSURU9YQjGezqRGl633TMYYnzfLC+Uigw7jAdgNSeV9eZj
4XkI5ktmuatFDo6f/mfZ/y3ArLb290RAzQ18DqNZR3lG0QK8L4zmrgG4mPKvyj4g4IxHYhPhWGKF
VDRHQi6hRJ4Perkyp/hKzMBDNzYTmfZaPQLY5bE1IAOIAqn7llDsChHYKh9HWw1gQwT/W5ysQ//m
N0fi9H5FqRX9V8XXLCMjaEHvLPwufJWKhJnReiYdo/nza4aSuCH0P2IB4xjEFDXAvREd5a7TJ968
GmjzkqH3/gCYploznwXJYmkjKPli7veHS8b0rS8kYnThJdaDiXjmcNDjhamPpSOe6MheBiQY6P+k
Yk4ws/9Rqw7vcRFaN5JxaKSXc9HCjLQWcBPWutS/uChc6b2l4KeNrotEjfI1BSVo4KQxIr2Z5C5s
LRlBmH796u0E/zLHtG6pQnNWNGLFngB/14kYrjLwhjgSaUZBBp5p/fByjl6s6cA7qR/jbDR6srwX
TZmqh+oBKcHd0LTVEpUxSoZqGBb+Cmx/tcVO5GcSkjwck1OKQpr69M7svFAAnggq5UzoAL/oByrm
PaX/7CBGzSPCs5Igrp315uBmtcauay4g047+Nn7BlqtBm7gS7GgC7RbqzhlWbmDBLY7W50PSy11w
X3KwJT5eCMXrb8wcnQZ7RCR6+adyizVZ7s8f1nrQT3CIpmMklEJN3oMi9WPujF0uC5jcOYGUU3sX
TNxOx2r48Kj6St8+xvr1QR+e58mISgjU2ysC/6r/Le0ffgOwq1ND8PzIbBMev3FQA2mYn9B4EKAg
UqjtpQ3YmkUx5R2BxLtlU6zD1AGU+BHo9Ru0k1VHizxrhT30Q5mvmbHCN6do9HR/ODDe80V5t5p5
uvPDRMQvAovxixARIHfvBxvZwYCEqpIDphXjMd4g06oVmQzw8SdOfVskxfGU9hkveH3Ir9dFRKoI
By9drrHBJ3ztGQft98SetmgM5aVnmECq2QmSdueUxcOcMQmoWkJUdGzmAnCIwE0i3ikB3wUeN2Mb
ks3b8tHwo7qH5Zmuc7c8HYQM7OyZAxU/za0vmrGEfWUZr+xYIhmWi1B97SRqM2DBHEUTfAfghOKp
1YhofgyIhAkaNbEA2DMP69qvbxkaqvA0PljXLijWK6K2pAqLJTDYbj6zdcHkTkJCyYdMpGsg3ZmS
jaBv0kkkRnEK1fMxsBji6jX7Ib23QLKot0V6ENus32nqKUvQ2h0ffhHE7YIrkQqX0PVH4vTMCsUM
U5Uy54mkQ2GdLMzYYJ9ocohIcO3xdg0iTH8THT+NGRKq1Pf4Zle1jnc5mLDaO6778IaXnDDWYi9d
K9NGcCEwhidhlS7+DCGY5oo0dcqnTTGnDU1zq3mRlglqnGCW3i5uwV6ofk8LO/KVdtWv/tPDKJcu
E+bwdxfvC2asgULbnFdEnhxiIPBHMjPmza8RTHFFi5QVj0rdf7XknDWSJNtO0GZm368Fgqmya204
gE7Ga6p9U/tWuafr2qxBAUQNPa3YpIbFs9bNbNOShcT3UQ/RSnhTd1HXFeNbFfPkfVB7LNTn/wU0
mQR6PR7OeYMHhSldmM/Uw8DZ/SdrERKTNXGpYYZBCgtun/K8CY25C/vb/tn/eyn7HA6SUNKbRF7J
P4xNwL8myQhbXo9VNpsUAnEpPoaN9G2KDXRmqREB6KzqYLDbMlWQ3Ddlrg3uRFxc6uKInk0Lot08
WhGuxSwCEehCHDFhXxVG02bnbcFVjEwB7KAMb2z8JidY8w9kYNTUMbeaAW8dSf0+y8I08rU2i+YY
PflBH5UCj2cgUXRKALRXfZkYhRCivR9pAFN2H1ji6UD8jpakFu/erLFUanjgiLxEcwrQ4uVVG2kL
A6emgQ64xOyaNvbNV+2EgIBDv/va7EG0saoM4L+RyAkrNvXjcEtCH2caxWY1lWOtieo6bZnQ+G1x
W064Eg8XfphGoJ0KbkXY5/pvSDx+I7EQdauJjjEjWibg+YjtNvKky4RSeiC7hHp8kQKVoSDMP8eb
m+j7EKTyKF3gSbFoqdzPc6n20oYkjLuNyXJ6ncmQDGV5IsvOgOZquSDzptKnuA84Ux1kpCxKf9Lv
bJpKsx97WURhR+hbrBx2T+MUAvPPc5+tysQefiNTSHD9lFPRsnRrFsb8AIHoYyyNcukuuBhz2q2W
T4qOdi1qLv8O2b68tXbV5frL2M3ZahG7weMQy5lxc0hKy3L1yzKBiK30nMnTFUVxB4k/N2Hc6bGI
DrHfwug40R4WpngMJJBYIIt7rgpMfoEJed4t1PSdt8cEDlJiVO1OBBx+3MXN/ZNY0hj4ADhtuyOk
nrzXP0ULlJq9Yytcz4XmUL7YtpV5zgPmobn4EjWD+0cEzXkrT/YUoV5MTlrp3FTSBWS4vT81sTdu
nSA9va7UVCPRuJ2nGtLCsGPEs1WbFbKLC7nDYahovkNyOj6KXuY8cbfceIxc+h0bUFPxRgXu1eF8
aaBoZx1fCXP11/9Z4Sh9IJOqBqhUOHb0d1SeMOAH7ZsKevO+c/e6xY7bodl/FnfX7PABYOqMk3BO
cZws9pkYCAKW+pGwViSN8Nhnh3M4Gl84/Zb/afl3lL/4BDF0EhHJxn7kQHHotH6rFu8iBK5NHORx
HgeSPN84028NDkLnjyOa5i9PrDwzmDhOfHw07bCe6LZvozilqRcmdy6PPBEGX0UNXjek8TszRPtW
L/5709uOMmiib7Ef5+P6bT4N0HfunkjLMTmbOoBKeDskVWQzS3BlpyYjqpswkPSEDlf3jlvFZVNX
MSSAHqTyK2VUnagpmlg5Mb2quwXrLv/ke6c8/C+216Uf7xedisb+YY64bL2F781Zok5xHQ51XPk6
GVnvgkSzYyEOSJlI0fP+twvwZrCaZ+TlpNgml2zAkV7S4OoElywl/XkfET2w22/cpEQlu9WwmquN
bobi6Cm+rE8imXhCYeS3+FEKFRgc/AxZa696wc29IYQSUYdTvnIoGVwkj+5fHJf6p+lAldvWYnqW
Qj1ASCRJof4kyW9fcdg4HF0HztJ7ai1IIvEFYXf1e19c9+/zyD0ns7Y8x/i3UBYmXROxgUb7FrzU
L6ms58Lb/H0xaIYsH0mJBxStmKw50oW+ucXZGBWrg+wp1dKLB7tWoFW1IaRXGfWLAj13FBdoovq3
e5OQ9hD70lIEwtSFLWr3u/g3ROgMOWDIwlSpUbLH0LSNSYlDAXAa1jBMoa6UaMWnxlSPPGHeMOvb
E2WfXGGdRg08KnLJnmWq3+UHT+HAiMXKN3cu8NLPmkc5ULVLsEdziX7PZy4pJ8hPCxo6fCWDZMYY
XaepGvqUsbE6U59HrH2yrps2X2/i4Bu5lcY/SqzAGsnl/fS8m7hFddvgrDOuIIAeeaRaNhnjK6MJ
oQgQY9s5hWiTGJeyBqQcqSCGtCI9eGk4+8yZqyy+ps608+qWVibUApj+tWlvgpTVwHJcAaPfaG1H
wfYhufV5HVqQt7Acf+BfEkzwzWgtar/B3yDiP4SC8f5QmjDHqsE7snHCrRUXlJDZ6n/C/bu0813O
uCml3JtqL+e4lxkxKmsClWfgFF7Uj5qLvxMwGv/hbFzCJFsmET6kcSQmiVUJDgughBxcWQ1aYlo0
vfoB4+ymfw/1Q0nqj8B0pgThNgOhgH1UXfmLZ1BNv8cUgjVWZIYZBCzCUcGeQ746JKCbys0JA36P
rhmnVNRgTe7wD443pjdCJ3yAmSGe8dqTIl6CFYMuI9G4/LTXRGD2MPVtwqLPauPHADIA7qIk4MA1
++C13WenjUwx5dSmVAhQhSwSZdCzflfiMmnubzmmkw0FjjWwpwXW0H6XviHk/6wmW6pIaj+3tjp/
WVOIC5rXZQxhPpd4LN8OAgWDLeZ07bLUBUHPVz6eriz/dgGicvVaEGqfNGeEC1EczU3HUn9dEXXw
mSJkVmja65MTYj2vdku15auykRu/DroxUitbbXkr0cFhb+91fzAPQ9YvWhaQ6yC1eqF2kc6dqj3B
ESPJPnh4KvHjmzzMVwpCsIWczIcQ+D9to1ezhLv4RHM4WCAnt3LWvsCzhpo14O5+pzCTLb6p3iEI
kdkxN61fZhpzUuTIsec6H1u0AXU0xfiVUHrsNVade4ILvyhTh1e025rPlIwaEA+ht3PFasnCWymn
5+p/jlR5P8Gl80O6dsEd6sRCeuETIn8HJqhY4wNgytU0zSu4FgCLQrRAhs+Iah3G7XflC2wRXbZn
6pg+7dVcbhvpcbcb+fjwtLKWAmfjS0nVFXpvDbYyx4ViU7tRS7SeKqx9w97hLbD8qsdmp3t6Ucnx
/++Qv+dzU9Wedj+Ro/PogrHbvYyTSEOpXOpMj9v8I52cv3D1JpnS8GJYFxqJTKLRmf/T5usEigDi
Pn0784RWYFg21909TpYnndlCL4CjZAr6j0p9X+yQN94GYtkXcwWxYwaPZqRmbow2yDM3sZ+AEOvQ
e01PloG5gkTtc3mwEAwKeNiVupjgDDuaglWdW57rJxqYdJJeBbQ6B9/Ku10xfALoXZlfx0IxHP14
z1ptZru+TkmXtnj8uCC+zCBnGRz3rn4gqSYP1Vy73EIkI8B7da+hgEFp3gcPYnYy8RCsz6PvXXPw
odwF+chZXqfSmjP8/TsOCcGuOZ74qpAgYx88nnc0IgF/D2B+wfwypx6e25jwjM4skNFzDsXu7GId
acufMcPbX1HI9Or8XmWt6ZOUO36pWA3hbvn7kU3xNWAsLtJ1AbyjQTIYoYB8QpkM4WhVwHd/bPx9
tJxCJmrFygSBdUZ/r7FeIUFoNgiHFMuzKOK9ajXoqvcnlI2i1ZS1d0yodbWxj67JqVfkwuXS46XO
szlGOzANMkxbMYmj5QCUWqVRiUE3+BQMKrfbOo9Uw7v+gduBiasf5AimxEenPTGB8QgXjBSNgfue
3Ao6iOhklrWzuxpbT77SZYCRZDCZaSl8hmei7KAsDBk+5aAcygVnJoYs76RJcx3G4R1vBm/skn9Z
6diVwQVFOtd/EdtaZZpSQbPm7+pQRk+jTxc255alwvqxV3LLLUnbi3GdCKKFsFWepekQXeH/g4h0
ShwQnqTkI9wRXZpGLGWGgtLl95I8Qqqxy+WjrPOIkrNrcgaemWTUrx7OkMVWMLD6wUhOUBaMCwn8
WxWdL4WglGa3RL7DwN//zR9giRb9dvWRLrfA1LEAZ1xvSmwqerKIhPE0PbeZvSW/R7a1R4AZJadM
kIBFVQh8uXe+eGzyma22nJTWCu2xfjykcq7/IrRpO7uOZljmV+F/9wSyUso2MdhlqhvUOrySITYb
Y/g/TbO+KCf4QfulESHJDqHVVvBfyAOjpMQxJW84T3RUcZqmOkKWdQsndKuR0rcas/c243qYMW1o
OttzX88tqDgxPDsqPi/M9iRrbc5omL1uemdB9jqT9Iyce/MOnLRxXdg8Frxt9SsqVyKcnFemolWo
+569Uxd7TpxRRvVQ56YwKbGPqMd5vjRLzCeaHIVXYhyj6L1jA/mJONrETQvnLiFCjY+SL5s1Njrw
hkWsrcIefP37jIGqEWx5h7PvgJcMyiWIY0rmorHEg/ax5bic/BtQYi3ISTUljluO7nbY3IxLxUdg
EZF0x9YAX5hQ/amqR5fWPQ4utAfK/g7p4YZJWmfMGAqJXRIQJQ52MmdLUA2h7sldRmj063zbPC/y
usESMquhZUfI6kU7IiZaSgASb0Sz7D43xNW7cDhCcBy2rOqC0KeMu9QpG4XbbiWtYj/kFZaIeL5G
OPIogmOGyNzQ2x0erjAY16KmRF/NGtzgrF9uxDPWBS0a0ewBFHgKSryJiWSCtbdiP4nhuKbUnbVy
h06pSZ57OgIq1iU70P4UTIbieZqN4UxRxj8W1/k88Z7fmrEFjc8bHrFyfm9Bmtb8CP5h5sIHNndf
qWTY5K1KImaDBTYQ1LIw9mcJr1bpHGABgOcUK/KNq6c/7fDPFVbHV7k4o8joxh7GeK7hbQwi7pxO
mCAe9i9LMfV1Bjhy8yRyj6kydijFxyd7SGJpxg6x6ZGtp2emCqaVoyAlGVuxBPNHsxyLjPQiJ8xh
BAkuVotaOUZdsyVvCavjmfgxO/YinzR7mn+dLrE1omT/2B3VIgfAf1oMC+EdweBmdNLwrdyHqoYB
KaVpJvqG1xO4LdDm0mIt8lJeXlx8gE2qi5zg/QtW+4UBc/LJLmBz1ILWKpQoGVYFbhmJXca7YaKm
LvQXDPfXgv40aV8MquAxygfuNV5ZRwl4fBSC/9sg0FjQDBjxQAnIQOvWYrMYEHPaU3woiINHRUDO
f4BjPNLS0wS7+qJQ6FQH+srXXMb3xIMvlqkneymRuuZoj0W9690ezHeMiu6A5KGI7Wj3f5eR6LzZ
WgSYlQAkQlnt3sq60kx+K+WbC+7dpwp5rneTTIo4bYrJj1ApQhfwqsVjRFrs38+4mXHXhxLuidet
hQDSbS2P5vKtnfaKZaZhDlONVvantApO6o5GFLNDKxs5uYF3lcdAO+tKgEKxOvjtjJ/f64ymZgHF
rFLdx5Yk/AS/cz14KSL75+93rhf4FCoFGcHz5AWyPwvxNHB22dPKBDC3knDNai9QRxkTjhONTvxj
V/gkrtst1+RiN9mHpAewNNrKl9r4IDyfOpdZ5GN3bscj1ali/GpkbHs8zTvOupdx4l0HV6KYVzJi
mG8FYyuS4mfeM+aNh6BtFuuV6QuZnO0Kfm7z0cuNFslG+/Nhgo6aOUr6Nm9e2ItFoc/jKcKZGpGC
+/LAxIQL7b/nWYcIfu4fhZbooa86ji007fKUIk/VWTeH7x914zHOuII2CtOaoWBQFpfWSPr7dIEV
rcQJJnzBnAMa1EUlPtErjVXcX8J7nD/1g+tN+Au4seqWNhnV7PaDAaSG9D3wV2P71yCaOe5B21TM
gAmIUOOON/6qdkLuK3stVXOESgMlG/QqT2wDJy6Qbi/0okRusowbPiQDtduXTes8zS6AJ6C2uvE6
p8YT7r6pua2KccTv8zAD/GWqEkNgiq4fnDsv5hHQ1yFITl5BEQ9FpyAJy1YlwUdlzg3H0IhyjKj7
Nh9NACsHG4c9z5xWB3y509ge9sKyXlMhEQ52DQC1UzA712q+Dgeg++mAFwSI7Xlr7h5dCOQ716YV
afWErFTEnmHyWfMurq10VV5eAKCmEJBpcq04MhK9Zd8HZQHk22sA2+zKz/Mvq1pdZw11Nfk3O6jO
mGAEcIvUJhQ5k9VE6mOF3GLG/WWe1UDiXGkSxW8p0IkUAV3rRT5MQQ1pVG74UEx/brPOQ3uqInmh
1yiOCMw1OgwnKNBrlmZ/dkzzsS+CoZ0/2wxfSzdzGxEd6gVz8+MYSDx3GOxxD7lS+gVmoUCBe2j6
f9Jgvh9aZFM2wr6fjEpSxnNDHvUnV8CcCXRhdxlaUNwB8qH9NMS+e6U7zAF9U0DvTqZCgsHF2Ftr
Q4MdstQ1nJp+0aHNNRcHumiQBibar7t3d3Pj78Lv0KaSg/xMfmQy+fWnlNGTh4lvR9auWGQx26qG
CuOYUe5YUzB9T+Tvl6koWPrRaNSrYP6G1x0d5m2e0EGA0o0adp38v4uuPGYZMclgtKk0OF+aBkYO
f1ug49VaBs7nYalsy8ZHShrVl1vKP8ijiCemoUEnBUSmLSIPgjxUC29LoNTmZlF1ckFp9qgaf+NX
NueJuOXT66HL5Wfm7NTFzW6nk9qpGlTLt9GDllO3rluz4duPw5xn0WCzWfsETfl4m1OMO+2zfSPZ
YuRV6h6LuE4UTRR1WV0wkKxSqU0hluYUCoaqN/7dU3G/t+h+8HqvdRjrPNh9rmuFlnwOKmti1ZVO
MSx4jfvXouYHB9zdnX+oHODFh9A9W8hldokto2CqJpjkvghEXQULXrgVFHLC3Hghcsp0hNbpANAT
joWZLfVgO+sopJsjAG14fTob25snOka1MRtCc1WeHd0/MIy1gTKCBfMkyCfegY2ZzetAvOzZfkm2
uvKMfFNy6QQq9wRuEW3OnDLSkPnU2Pk7KRFTAvhExgj966B035/fEFO/oncU5wjM5fdUeCYj3FTU
Uxh1ZwM7xlvinN/eaObmApRH/z5IbwsL5RT2IWH96+MkBQIJu9jAb/P5LAHOHFq3T0VNybNZVHhq
ZBDzMqzjEvVIShoaRFGLpHA6MRc4UPd0ANT4I6/WFdYmJ38uwL52sZM9P6bTf5AS0hHAEiJDpV3c
P883MNOxtraMUAO2nyEXSBiemXY480BexYtwmgQkNPEwh5v8yyoXGbm4igSUsACCtaLEr9Orw5Ei
mbmTzfuEM9iyheL13CABG6kOGUW1fLtFico6yakZBVOrHgaXc5V4oQRinYd+0weyvfi+Y0dUsBKa
mGsp+xODs3Oy22hZsI1Uqypt/ixrZiQJnwk7lApUIpbx4/BoBEqd9GbcHut4753gCOyI/WFBnjS8
OH9/ochRn1ZyAzdEsO4HfUZ6sJQ04yuoE3wsAIWotq4h5s4TuheSM5nfp92MyLZ2039U6NBMnEEU
TYEpc7OdFprQpnc6QO1IAT8ASbuzxGoN6HdNdqYs30D1REIIsIPYXuKqx8PebVFPd5YAHT7Ikxpa
QArScQ0+wkLUsYuUkUWCY4h9bi3gxR/5R+ANxTFqSefcqCbfKN0Cqr4w3G9MijNM9GMnDWKzpE0s
IyfrGT/aLUTgKB7aUzIsqmjfQmB7BrsrVW9lBDW3iO55Ng9+SmzzuDWj77JZHw99DRK4Z78VAqsG
bg7c4QPnlUFgip5wlaIqvXtg8isTVs4hzPaE2ym4ZIxLHDssgoUUs3FCtZJbsQP7nb9PG63fYg9u
oRd9bwDnyUm2CoX/9x7TUKuUGYskpWEj+lRIK06arotHCsL5fSQCNSd9kM3Ahgq2/NJiS7BOZJb8
Zm2uqNY1EwDB1zQ62mr28A5vP62bznOtSXQXgQ796/SqJ1swbmB78i8gWnlyPLATgk100xu6aMnl
TjV8sZlgNtwNnywIQUJrktx4f7hUd8j+zUhh329Ne0weugXCXLsOywxAujFyQwBKTgPBadqugjBM
UErXcA8ghhDUO+9hJdIQR7hb2rqH5/1lXq3O7V3waCuEFPGqcsH6wlUSC82hx1oFqJdFUzYce8TH
X2ZPhQVHv1ZMZaQfyg7nvbhc4f6Yf0BVVIf3UbIEjqID+7GFEg+4cM51PKtH1/pUYFOAs53Kv4I7
rO1r4wAErQU7RnxbOwU7TcxxILK4Mh7HQk+gWCaPB7d0aye9IjeD7yTUtoEZoNW/5pR7WBKkXlrF
NrxYBgYLJKjDDi3H924NLGSIQploWYaSs0y0fbi254iw73YLHx3a+8cebz4WXh2zoTVbmhzpeFks
Ba26hRNlGJXsXJlKYqasLenn12WjgBfkos1x3+OcRSls8QEBgT0VIVaJHlbrkYUeMyEtJF7GX3n2
xeRVZZ3Oo+uMd0U5BBT2YD/AzsopenBSBmEDR2HMNVBBNQh/KhHfx0Um5QdLKsVCtOm3r3WkvQmX
T3/O5ZAKsvi/6N0Ibhbi4f92ylvXt+yAtVIabMj8ex+M3C11Gff/9d300e7EcnMq1m0gwl4qFyx9
fJGyHR5uTwaaCd+2EYOJpgxarZyie76gPjwlIaIzMxq3jFMtcAcJOpvxMMq1s+36I/J/c+4nR45+
tFsMPb303N9ugLkIxfkZ0t+MGih05wK6HOycIUSd8/d7Yj/fBCu7VW95ArE/zSIXor+XBpsRqwPB
rmu2XaczH5+ZsmJlhvBwuoTshR72+HByKkFOCNqqXIwJeod217TnCkoJbwKv0V0Xkr1gnBPx7SEl
zyHyU0KOh9g0CSVRCITcq+coKwvo11XujQQvzX35DhmiUNuv3/esBD8XI6J+6K8o4q3wGA29C5QH
DwwucEfpLtcq62WHnUwaf2DXM1STZEe5xHhEHD1XXnRPflsNNL1BP7UD4Ctor7sVk+syLRcY1Uj/
iznEwjrCCYSVUtnoync+oWMhI+NcVHXvaQd+tpAwMR0xzQaVr4TM2/Ho9XBHhFu9pT90MIKFKE0G
NpmnEKu4MfJFFReTnFZmKA2qnLvljzDZPA0cHlahqE3LntmsFMOg977k2NMxzgs8WznhB6ge1cBf
kAyaF5T5RFbFTSnaXRDjYkY4TCjS1kvEBrA6c5s1VA3oCWo6LUJUXzgvnRpYIqoXqXPOvPMt6G9f
cCYMhOd1OvlwRNOO1Bctbk5UqcGNSuNHdk7Iq6tPNRwUSoYqHDD+I3vZU5fGzpS/FmdPZGWKGrSu
3lIG/KFXn/5zJCHrgvvpjBa4DK15Zq2+4mzvq+mH8qs5lf2R9PIMaiM0JXrnnnmFc2jXH+rlMU21
QZTb70mLF/RYxTS++fcq6CjpZ14gq6FUdTmNZ7pxfh3ul4FgSe/CGo5/Z3IAnBM+XZHTDElCF6aP
2GypHVuj5KAwXmBubGccPyP9kSSkjF7WkN+VBuAw+19/WizGpagSTZxJ+UcScygkjoUqOZYA1mZv
Xt6ljWrcu3Q5gx8KBq5+myj/KHO4zuwxI4fZC7YxSa4EtvZ3nOcQBExiFgDaOQalsuqtVDqOn/sh
JRWYvTJTeh5oXgS9FdytqAR/w4tcwUdiBIT3oIIL4pEzO8OHfChadvB0y58Dl8CW97VBjWA+/Q1M
Zq2Vp6XIkHWwPkNTM56wVCP4nU5+rsHRO2cwmLwnvnO6cnRwNthMWVBqdohhNPF7Bs9lnVUAZdS2
qMQngY/TCs7wQgxV7YuFK3J45eH2O4vtioQ4i5BNJlSONBxFFV2gXRNdmBIBGeWs77ZoOYqnc73z
AwMxcxy0Elbuh2A1bKA25x+qoQmuRBw+3zw9yMTi0SXjmDr0mHm36YrPfFS1Oz02RmrAInf0BgWW
LSKfRIaStp/hsmZvOlmMSpwuNyWd8OyBk5OJYJnI7EsqFKV+Z3Qxe1mXy76eQYRdzEORU5OIkEB2
fpzqTomBkDiEut12ZuqP3775ia8XM1f+iNUnOy1/EoDoMmkNMpnK6hhJac3SY4LX2TX02aDgRdOO
3fh0Y0zGNkSsGMOlsU3YkYhpjQiMZTk/YY9s5vSB1H3SHk7aP8qZ2qBqHyhCZDsvM5E8kMexJKPh
j94UT7cGbWy8bs8gI81x57dOGoyB9IwuovoagoMS07COBYu9o8gH1OrSlWLkBjt8HOMYkbQdNZAZ
Du4fRSAFtFp0cPknMH2q6XjeUkvcphYmdrUYMmMH7niPx2zEHdK2jVohup/c0k/+cWXIbOzTbDZf
Xnx82hBOWiHaGlX+1FSMsqOLI3DXOABmzsfcsVbOO3wwJGnyA/yXq9F2WDefJXc/hOV30w6/VhD3
riYteHTb1iyhO7cJg/FwLtqLJbmJjoN0oYK0ZCuxIaISoqEHOJtj0HuCDHC32yY409HiGmURdWSQ
PBMZM/LEOqYejMwJofj1kgv7Wth5csTPlCkUt3AhlPo4JLkidOYb2kKa+Sya5n9lT0iUsvZ9t/mv
Ly+XdTnwKp0tswqo6tYQE1JNeFH9h8UyLjZ1Gj2p0xwV/N/DJK8n+juvQ1pTxjqgoax77u0MOi/k
d4vaEo2xhTDAJgqXTmhTC7DjirnlcT6zkNZnkBbCEalqksVA0D9Z9/t2HxcmkMqBvdwwRSYQcflH
KTd4r/7DlnOJqz+Lp8CI7UfnJvHvtOg7iWADigMMnURgOfXTCKUYb7uqJv7I+p1TK6RTxB6Frenx
lA5l+pRCVi5LQgAm3nYvd3DdOAlZMM6iVutN0TtSHVGPR1unwr/dwNUa4bh6TVy8Wj44iPmGS1uC
giQqITX0IPbsuB9n42Tg8fMBwHetGTn01xREAc//ylyxwnFksoct9OklQ9zNJg/W1dY2rlusbcqo
CqJvpJNiZWd8ARUcM4/cZrl6LNy6MhQsXAkUEwZsGLWRPpUcaUr/KYUDh64KQdvz8mMx8dHZSxnh
39N+wMd6zDc90sNlmGwr/4Q1RJhy/6XhN0RPFO6ngzzditJtHwWENayam8s9x6Ku5PReE9li1rGI
yQHEEA4lqsXcvqwj3Lxy4vZGPEpXkOXfbft1atne1W+oR2Y2VtYgfSnrkWdU7as/4iniAvn98VT5
PxiUiNLoXBBStN9QteyOdjhircrTqqetrdbcXdAy9c59aSLu6Nw5xxQHX4c1o++r4Jflj88YO/Fp
UyrYaScqM6uAl+HitdDPHNvCWG0ZBHVgcrf4a8QUJO0YLITMZz5ti0kQ7oA+5unnHXdgU+mTbEA/
XBGHMXfdFvOnRd7sHrIBHM1/gDVmHmbRvs+BW9Sat/PQkKGP0IvWgt2JmThPura9LvCGS7FwvMCa
jldVQOVuo9HBDyBRwg4wSDxTkwh3g9vNG+YkemYR8dMBBWl/Bw/JarpF5Be/7DZ9MBn2oahgzqzm
Qrii2au60EppfYlsXe8rVFa0MHg6ms4/ituLtyv5a9kYX8fBTUPTEbSV82/hnx+GXZAA29xuXXgb
URHu7KiFO4brUQHShYY2HxH3jp+Vq3KZmuMmj6ToETndD0ogrgyN2SroTaT5LDqCfMjzyqM1Ll0p
RMo7B4fCI/fMT8e1KglznS9p7XwTft3RN7a8wXGS1uNtSjJGvQpP4hKov/qZNTo0lM6oiPLHKlcD
uNDBd06NCkAXx5qhFljP5sQOhgn1uCz0XsCWV/x3DISKRsLDg/FFJoc4chSadiconC1CfneJiQe5
6rfPK/G939/vl3SxDMOtCmJi9EystJK9FB4grVe+ANS7zc72BFLRy9Re0VNwPStOaY9uSIw9TVbF
7V0UG2Sh47xu7JUVSwCEb6POad9RmMmTvH7RAHY9qcpDDOiUf1K2NUXrU3hb9tcW/fWTjiKeaMty
48s2sTgHC/CRG3CzFldqYzbYBl+JDfGSNvRjrEZuRgNfeTX1V1GjKZ2OUIPLLWygJe+JBM2XrqMv
rxYSNGmAOHIpbs+++22kPRUb/Y+JghSxuCWFZzKLP36p0lhwBkJRSgxzmWvhLFSzIGnSTGVfBBpC
46NWA6ySSCQ/jrs/QnbUR7XfAkOjEIeUjHvNgOYDcozkX5MTvcmcw+ENb3cZwyV8YK6tG8F2jNC5
UntWyhtIdrnq/4vNYfYM8Cb+bqXlVaVu52OH7hEfQZUblqYswyNhwMqv5AH262TybMfeIWWRpuUz
xr8O5wr2Dh/wd/AmW0Q4dOFda9yZ4WGO0BaIlTVuIUMjjhjgGzQTn9Wyf3zuxLoFLVZBLXSUj32m
YcgkT/yBxck7E/CUGGwsU5zZJl2kTeX+jmw9VkjjWlmkVzcMtlEUF6MaQ13az5cQ0/fzgjMlZIb6
UKlyeY7O98IpIx9YL2ucoDjME/R4zLo/L5gPV2NsA5V9BRgcF4wFU5w8m42KOKpTiCmsKZ5vr+s1
a8IH9P/O3IpeGmBcCZkMWdPvGJVlDc0dEkgpZ49ATs8vmvAlCMZBWATL1H5L2xK24dNwX1kdWYeH
mCHKGS5ZGoJOsZj4RPs3mURrQX2AWBOnHWvkw6tfqG3KRPOclAPmSVrPvpQW6lwCWo8ApbiFZoav
jyo/NatGhqjDH+dsnqdr/wUZmNcYviHf9/PCSqtRzjEcPPfpTsoIVgGCJhMXWIXrFM1guX8EOrAm
X9mhGpVfSfl3dUAtn7y1qXAnNczKcdweM2Hk8v1y3jq6/ElxCfda5IBtRwE4o7oShmZ9vea8GqiP
Zf7D7Ds+wXUirPcYLlpK4zz8pCMKtflJdhNiGh1a7HbCsgX0jIyl5taYgae99rKJXhkRmmWbMQk3
yzcaqGxEWyt/SzsVQX9IFQEHx1QdUsLY7YtK0oDSBOOzyqDZMOpEKAXHYZkJr6jiaIJmdB6xdsOw
ZWON4aW2ZmOIrEImi6Z3zWxsgzzy/U1AqJIQqTX9WBZAiUsBCdoVG85a/Tf/rrKiXkCAAdm6YXVv
uZ9IN7LFYqCLSJR9cOzhC8jTGq2Ukf/xguUvqtfjQSlJe3X4GSNJX2q92XpU+hOYSfHE1uVxngL+
B4cdetIQXbPeciSHXkrxsyEOO+OLbSmx8LTEGCWDw3oIEkkIBH9rG63pOfOKYWTJ5Vgc7Gh/LHS6
NB13JWai8X5o+9kwrVnJOcH3+o2ztffskspYgGkHgcabOEFCPmxYS+MltPNK1Jd/dFr6Dq+b7FKR
j32qrRj+bIuMHI+Uud5StRVmAdaj6C9Znnzkhz/6qcmo2Uvfzt9WS3EUjtFR3/1+6qoK2QiBPX/F
awiK+H/6+nqqfmEppbslh3sO4f/4yO4S6E/qU/m+sWfangOlCz/gXw9rfNzfoRBNkOnitin+d6eA
dG4ubOtrYw1x+dkke6K4Vz8xQeMG9Mb/N+hyXdtPFgxxmO5p4Nkk4OmrWppu1B/vtmkphTAsA9JC
GgKJ3E/TDwIgGTawhF1A7FX6/5kpo8o2DwZGvzH63X7gQ2/Yru+BodCfuBEsc3PjZpMWcpYbly8C
yECgOv9q0cY8mwuSXaDTrx5y+X4HduBUT5sojnZWKWSe2MWtaGF57O9c1XZgVC7K2ujluqDvu/Oi
m1HNRiOExraqP6LrW6rnrRLgNwm9P1qbAXVB/IQwTJzHf4QcLYAmgCfSbl3Mvt0ZXNiNgw0CUptS
49zc/2HO+lvRnt+V3lUNPpvEgKxcarmmyjs6aAtBfMkd6UDKRO0LzRGmZDyJMHI4RwBWQQ/2cdCN
ypBuAaaxg2hkEuQxwckHimTqtm7GpYoL9LjtMRxqo9LRl2cWK62sK20lnniR6y82+yI8tK1QkU7z
Sq0UE0I0iTE7oqMfml50KXv904y8wN/tQgAuEUzPJPT96dV5nLHVaYRmkDjGDdWzGqfYkHtyUVZ/
YO1d4tq6MD4o9YlBMSg8Ud4xwoALTx1Lwo0ldKlL73+DoTCm6jwO3C4BBgm5xn+LquDA66TejLK7
JsRWaLQbEIOKIzR2TZNoWtY4PfYpYA8VdnfOw+IuzAkFQBtayfD6PTyUJANbPm1TvjIrixlAR19y
Oob1phupXzCrNqvlvp77W/PUvTN0qO8RKm6ueBka0FCU5j4G57Jw5I8G6lekBO+J74XMAD7u/RwF
1+6aCXTw5Si3dzh07z5gwawbB/LWarKPLz8L/x31l5Nr6MIDrfUq0c4HIRu7RX45ng4Al/pApxyi
DisWTc1C9OaOyge5bdc39ENhaiUit0knX3f9IfBGScCc0rCKB+jbsmpLnWMeEtTIoMZXxrCL96Yv
PUGRFfWLrEyQhfXbOXgNKzTX0dFCyWnuRuKxQlvicoG/DS8Hrp0NoVF30mMWIRLKoKYp+OUAiVo0
VFoVoSnWLT+rjNwJvT0JlZXNrmwFVuqT4Zt27Eq2xr1M5XaU6GhrWebIJ87KPnlO9fP2GawTxJHK
BNKCy+sQU+C0XpYqB51hGdizGCg19AGCRmnNN84Zpt7qMlvTwHwi6IjG2hFXyVEiYhI+7CYBTrYm
nZxJdtIU95iodwAuJ9qZJ9tsjf6wt8y4cXCJ9H7UTsBgL9JDjD3kreSXGG96yLZEKdLFPG5U+jPN
YgCl8WlXnx6HLHgrJcH0eIujuuXEcUzAl/fJe6no+pUmrYrdL7RVb7vQbOTTZqJtIUo8vhKe+QVV
FMXJZuW091IPynQ3/KuxnJ9tKNiwltJwbMkZR0bFiywTTUWyUB1FsiSwhHBNyvyHpZRzZoU9INWR
hTiraWMc5iwqhUr01l3ExdNbiD0gDB29fRSmrS0szRT2kJ+S32oYsyMjMjpFG84zG98bAqrueoJq
3mc1dr/vxeuhH1am6x/bQisJTuPRqFR9ND9h1cc4rP+d3ShzWYD0myVAZiTxitcyv2L1uoMarBI7
0iQRXLlS7LEEnsfRMzoCpoFcVAjAFdndGXvCBwCByzb0SZxHYn4Zn8ETeE6+D7LhpgjUuIPMcI5f
XdppNFV5DhEzeO0snkn1NVIclhUGRKkSelP2TNAEbdsvNrxpjSzZ5ML9mp6Qehn6CC/7XB5sE+r5
8Tjr32L5DXlbGWgAKQkfIQQFeV3vQULRfaifgb+1umpfIAVEIWS5kxVbuCObopQgDxbQep130z49
x/sVrMntmKE4q29uvnIhDQ/wEUNX1FOtHg7ZQWQiXx/JuEj2gLTAU/kSQNUstawQXklBxpw6Z6WT
+bM/lQwrNOh/9Af6VRQ4Xf/QRR1K+ao6/gpTiQ61s/+rYDXpOw0qqSJMnG4RGP+P6DZicmudBeMC
OAQfFWsSBFBwHCrl2jwS4E8qg7ux22SommUB9A8k840fd5sJABKv0gacM2xE3Tv5waw4tvM8l55D
lt2vC5Ee52hfuX+8fcAG5JQ157+IfVBZG7EUzXAsyfevH+yNWFEQfWQU8gcDqYZ9oevqmqYM8ES4
N9CBbyoTBrNqXLQN552QpcXC3ycjzBkGX4IiBZ5xoez36y9R0XVUS59bf818Kg00tdwJrAOS/dd/
anQLFyOYRQMa6bWs3RVzUEJhT4BmspnIEnW5srOT93r1N4YOHIyWl5yz1hcfD4bqC2MqYNSgNoVG
EixCgnBB7fbMGIIpLhxH3QT+xmjC0Pb25RtdJ9P1LOKmXzcL5KiMVzvc/SoOhCUwY2iCxV7N9+mg
j/WwlcQsnEc/UP4LuwO1shkTW/m23frXsGXjpj2yx3nj9JHLYWQS5FrTplWE6vS6pBfqdQDLRdeR
+M0fJzdxyfk7/J2ErCpPLNtltkKb8LD5S7jlryqhqNnvE+vCRz5OhSHqfGR3SLAhnhBpalJCgdyJ
8GGu6qN5Zz1rDCUUfWW5hY1tPDNj3jQsIsSj7Qy6BSoKRvGG5pollsu8kXdzq6ihqfW1AjeFtT5F
XRyG7ExsuGcS6xN0n8NfkG2V8aHO0a8ep0vlRP0GswQcNPSvMgCuHEwmtenos6Jz7AqLjrtMwrUD
y1CI5bWCTxvni8JD5m0Dpv63UBbiD85G2XAwdbI81pcby9FN7PmXMh5Bb3zatS1opHo2sB1sRy0T
wavThAfV4k4EaS9PQPvl6PZ1LqNWtEfFPWblUqNAurvoV0CdtrqRXnEo2v9ZsH3W/Alft1HjM2l7
wy32xkYblLIqdhW/KDRv7qKlIFeMRfeZx9pwnRUs9mVZTistjJG4VGyhrID52wlpceKFna51m4TM
psZT3BBXjPo5ijjFO7utjWJvJxbQ99cExJOGjwaeBmVarGvAmKwqhvgfXd9Q7gWVCxJFwbJmbvvP
GgTVvZGVuCcvxbOT0qVG2HatFDQAGf5uHjfYYrAGfkKHf6lxVN01PBp7Oh8yZN+JFpnWXov27Lo0
k/XfMfWnUgwQC6828GNfDKiJPWw6N4TxtJFlTG4VyL1wwm8ZgQRvsqVtVbBKnUjcPvCxvvKMi1Cr
Mb7Seia/TaihlwCpXBftiOlJWGTwOIspCZPrUawqW1FoXNpoqKS2VoE/gHCPctMaQsalE0MaPxWG
4qWaDVLmTi9dzDQQQW95Ucy2wKLP2LIwntGcksk7mOWtwvyNFJBmQPK9SLSo/ZdswIQrFmqGgosH
YTM5Xo0CmeEmXSRQNewMCCsBmdBu4rqIWRymg5SPmGhCEJqlpfuVXYtOxwRKH/7BiiTj8I4BV5h0
WE53kStbH/iBgfMm3cCVjUTffecyC7W0BMEB6yNrMbWrMDX8h4JG5E6fEbtYQ/ediGdsjTU3yfXx
V8s2cj0NQYo43QRNJHziGnw+HODBjZf5utZ8DJO5shCx2w64TrZMeVX+wyabvziDw5XsUHKUcbgs
i+ArrSyFHc/7jxTofwQco9bbZyt7AOlWvRmPuxfsIP0/q2LUtP3Nzmxcb5SXhd2YRSSCXb57eouS
EcW2ZdWUffrvMcOVumywD+aq2SrA3U2xP+Ksz8yruVOb1LfP5Yg/ugnpDDCOq50A7b3tWd5gc9b2
4jKjwPwJmrmqi6kYJUtJ1lSma0WRGudPbqhPtQcVNm/8Uxa/rwl9mW1fIpqw1gcuov6FOIe+OF6z
hn5jfkqOa4Z6gPxnRdxc0noybzJuN5fRSEtH3MW5BuhwQpDkyu8+dDOh+ma/WlKNCPbueS6ffJzP
o8xzP3cXmZKFwWcBHl7grJEir7jneoeNBMPOhWTCozkVm48RjzZtdoK/uIGM1V0s1AP5lc9OTqmU
yJaJ6mmfCyXhNSpm6KM+I2z9xL7IfN8YLUe2fbK27q83/R7OWTYGksGA5B3UKOJ05r6LAEXFvF+D
YsGBo3o2cGpgqXjD6Hyt4hk/cVKCfZpy1iRZmMOYBQ8MDV8g3tq260W1CRIdvy6n667YN1JTc3iy
YCAEVqFjFetao7dRzKgXdpAa38GGcptEgLWxaXR1QK5S7+mPp9KhLVcpPEehswdLQ9dGeZ4ReWf9
Y2h4BSpRdi4H1ouXsSw1m09/LCiELIgsyh2/b5ZZGhtd+oo17ASOZXEiCgOTXuwYplRQVnTZX8Fo
BrzQJHkrZMxKcc30Hyw0zpbbeqFvOR8yAI26H7WbIui+7DADEt1rGsgIW91bTVR29mlRgV40ZEIl
/3b353aG2texM+i7cUCNURDCydGcLb30PwCR0YXfFFIt5mat5hrLx7evu9yZ5SQ2MmzdB5cg0DId
kyg30xUIejuUJObBENV3or0KPzHiNxc7HCv6nioc0fMVdRqs7S3UkeKbqQ3vumU3XvXtd9xiqBZ9
GuZ1HQk6OSp9f6nyPl1CcN8hCtd8jL+H97c1leUMsh2i49eXmkxDy4XhUjFSqogfgGXhJ2+fbtxu
223/hfmVe7QTruIbvpdHKsOWkjQzUIoRIkclldf9jXxS6OjPHuu1/1INsqSnlT8mRgwCbFLN0dfO
Pl7By0j9x3+JejPfVmwngXXQg+Ig1p7szZFwkQUfQqkYBxYCvHWvJDJweqQBfBCybNUikUAuLV6o
uh8WFi2R2n2EhyJd278qDLKZnBEGCl8wf50DBLiy+v22rRZYD8Wsv2ifw8MwsveSWh+UhFR4Uc64
ZHsKYNUryxXjTkq9kkRRPRdAayiOpaC4mhVj6BGZ2cQZZYh9eNISeagpZNcA6ldixjM/SApmwTcx
TYPGfvIdhH/PiCesKEy6PrAyGLptlxKPc5gJOJso66e3EVsZPWJ27SGlGdemBSiFyPZFsnc6Ab7M
ruj4v2XOydcXuy54OiX1EQTejx4bDpJxxPKW8eY05axGGwOEItiCXySVTQbtUu/h8Pm+XZKP5YE0
QGxEgNpRK7vud+Tc+EMHCdFOznvm4JEFsjimZlCctDlIt8SMXWI4sYA7BTrSZAj8MwoiVe13pPlC
23UxmIQuzj+mPfd8on2jLcs2PzyhXrV1wkV4ngoIiriqzG/PNQFwF1//H3P9KBZajKniQ1joZvzf
aDW/LJZFgD5j69erWdN3/Owxxzxvv0ApmdaQIr6llMxqvG1HpZ9qJSIrKOevw+Ql6bfejZQMe4b1
E8EvH/7TGexUWb5REg00QsHYcAv0gipn5TfoHJ2z5lII3IeRP5iRCGywzu0CVZSA0mxsYe3BDw06
H/U4F6yvUC2LImoIAGSsK9BiifKMRWekwMs4voZrC6EcaBxxK/7VU8CT9KTnau7YYiKUCc/HrusT
GVXPB9FjNYZuTKzTE8XC/36SyL0qXo/otpM2SRiXfvSoH0NpAjGRKItQpY3OL+pX2KuAlRCABWjt
l56aiOGiezTlIsXm/aTX4uf3pRISBFMYe2VqJIlOb0iAi8Y1KgfdXYQw92Gk6GnaPGJQxCWqGrNA
UaVMBUVL6jAbi/AtWziDI+VagpaI08Vaen6qZs2MxbjTRiRliki9UrQX++uk3mnZv9SgIxBevo6x
dIQDcc/V3jX4qBVsM8oj5d3pkf/G7+tU0cFydMY1zs9Im40V440LnJK+Q0e++ITLbsjPMlSN7Jm2
qu9Y1C52mVsO4qBpLZP1/9bYb10E+ooqvZHDRrAHzXb1W9ohjx4rGXqcu1bNrChQuCqsxmiw1+ww
+7dO5qbThfN6W/hK2duNMVEMS57SXA6J88N7FB/0O3k7Bh17CSJ7VPfCDG6bhGHddkQW8g8IY10i
pY6tz6XMJlLtHBO+2Rd2KE8WYIS3Tc3SrlaVtaMRZeWu+qT5SRCLZdYEqCceXkeGVWjr/e+LL30X
KyBrweESUDvHIRSVDwEcPCgBFblky87Z1VVW+msQ/BGasQ5nULSuxnLFKhSGHdgFuWGlyRrPlw8C
Hd1fkG+UBCBXZnyXtNhe3O2rC461IvtdCQxkLAJ0Ts5ThiOleXMXaZzA1cWIpu6rAx63DraAAsRB
MMY2CU4fbcLofVkS4ZRqCnFrx8d7lRt1bWp5p30wK/Qkwz+ELYDQ5EjPtvMfLktrehUu0muDimVj
EVnfNDOzKW1X4w7mG7csyKmn5Lf5nQDQJHyWMKUb2tME6OzEYUVDB1Z5ZYYXwj7qwJU3a+am8lI2
kv6BM3g/ZeoRZtCR5nU0ygIVpWZqfLZqiDQwh8vO21QmbcJkij0P5uyNQgaWq6HRii5xbXcWEnC8
F00qtJTZOJi+K2K5u0rXv+92NYry/AS0TUh0kueyErNQBdf7bu2PkBj7xEQOnD7dBZUsD1mpiwzi
GNkcZmcJZC6u+g4XXxXLuZv9lZpfvUbyibjdxYNycDMvQ9j08bDg7XDdK0gXNa1sGYXrcfdfAtxX
++fL4soblpmJIEBE0yX+QGOuW8k9ltBWH7TlBm1oCie1oQ8yf46whqBKoFvF5fjh54+2bEwjNyk5
VuQioObAV0ZuEm/PMpMCMObNecUhjLweyVoVgS4VL1oYZfpJhTxE6K8pEJCQpTjySzrBk7NE0Exe
sMYme+RrbU/CbMICTn7rXTI5gGGlyvpuGfyIDIlHCNhkwVReTgIWSD7gXoNXXlH/q8QzenZ/rPF+
3YT10W1Kly4NjiEDYY4LWW3JMuswFTa0uKI0jbAxqXeC78kU+8HMWFPPa9xr+dG7xJlIvCM8qFxQ
0FsxB1VIGDDKQfEq9olHaVTsX2CCq2m0+DNl1oedRXHlI06uQrAf8UudnjBh86k3jrf+Rn/QLtJJ
bUz4IrzDTx9R/1gPxLi7g/97cmO5rTOHrGzSj+o327FMN47ZSODebgLsw8iTmfjDMAQR4gA2PFJ/
L+oWQrVhZk+PmA9GrDsbt4/2xFGKotoaB59jBMhlWjiclxenEpBZ8afs+blePIHZYKBqLDPRuKdT
OCwtxJ93rrtFrfNpdnJknL51lZu8Fgu4/JkjaxTYp4c4bv0PPS8f3cd2N+d5QridS+2QiGTayoUa
b/fFrsubD1z9846KBNsugjb2rKKFcDvKMz0e5FnYv2Xz00YlNSlM9zWkxpd1BkS9B0HvpTBj1mGW
qZ6wTu9wV/EsDarLoxnPMZRZ+ALrCX7VexRix8RK8LPjE5uezp+gaUDqBc/idBGHDYjSQ+nfc4G3
R4okf8bOEGsMaiNUMeybeOrTcGMEJxGw0GmuuPx4wEk7xDZRZyK7OTjwgq8Ya/mEU8VGDgZaC43u
PSVPUiWHe1DF78DturOkBnCyQ3qtBHhm1swyV2WW1Solh8QNpfH4NYYvIs2j+7GzBvUsVKOQ9a3r
FpqL+1nj4XSZats2ji/1ztH0Ym4mn5RU382z5GePZkdoHdoWVqEWo820qPDme5cUCrWn3sXIwf1s
K15qvboTDd4pj7PlPXvaP0fCVbn+iPBMGAOE72gbMU9FbZcJsya+c7ZGe5ztdYkfJp7/1nsjOQkI
11RMndvxpud+n2Fq8+Yc/+AVxQQki2c1dDXx0GE4QDZfPyL4xeAtrCutB4W0GijnH0jQPAiYAMYM
AxcjjqQM2ViBWCJlAdOmZ+OFw4Y0fRUAWwr53FcR1AEU2bkyqh17UJj7WG3J8jDMpt4Q5AYeo1FM
voOlwwiMSZDIlsYd0BsWg+OifN7Bzu5pk2Kdm6T1ABzMn2VSe+EKlAq+nbJZctMgQf1NZWT0DIEY
YQFA5VGI1pc6Bc6OjrkwSZExFz8NruNGAK6ExzhrTpmAIraATL1PoA3AZ9txns+hT6XduJeJe7vF
bq2gYudFov0vGpLiv7XG6H9cytRHtw8hwZRgWD0NEc1Yu9Hg4ZqVGPABAG7MMX/waRfMF6wX8yGU
O04kJIBz54pVm8krI0uCjVgnRe5IKDGj0LlerhIcFruPW7Vl8ba+kZvw/96ojWG9BhVcJ8QOF0bu
yW9YQkkN5Fzk/38D3dblrfgPzWH8ByqrOQ7/luR+A1AcMS6MEzomLxGMWQ9F0pQULmMcELXScpSK
qJzLd/NMSIWlZrJIOIKN9HALcR5OtlP0USrfPq71jTfNGh13KG6Hh3gU6iu1ol92mbPrTTrdkzsu
xnQzl+89u5kbD69uFgqAlO9LLr7qax1ieN7TQjvwh6IlBtYQWOD6CiY/vt5EKJs6wpMnXUpullhJ
TKcRF7Fv2Nl/K1GT6uB/Vdf6lU32yrBn0hcSj6Aia97Rhn3B3sjZzYMz02vprwhMeOTJOAWFBScO
PAOyJjqDqYoww5ksHSedY8eHfkxBW5lvPumdzfoHn7V84/OU3loNDT4GbF/VNa3b4S5CLlm2sX0t
U44I5FYqMF82YmRA6rhWcgi3kqJpp97bIJ9vOFnfiI3TzYthZ/UcWPJEMZfrw/bsHrAOlBqetZo+
5wbw+ndEcAZ1hd8tFvgf3nZqp0tgTGhuE2U/ID2vEDcCrH96frmlLW7OjG2Y8VAsEunilobPW3v/
6yglhKUzCdUxTjrvCXb7WbFhEiZgB+ov+pqeZlhLBmeoO2eeO0p0KMWmfAiW48zxUeb58d70uYRK
pvYa9W2jVHcOuBr8DrO+GUAuF431/0/mIpMqS+8GzWQVP3kmYQn2X7tFnE0lBJw61ysrdbWSxE28
mLnJJQwotiZrWpbsoPpVfMjZOV4+eDWLBdOBqAEYlaYu8VPkbvQ9U1/sKGxI7LxKz8trTJyszLnM
WlZzI6BslkoA1KpovGjnhOK58tEWVQXnWgT6Kab2vCJqzwHa7vyMubV2S8H+BMN7+DVQ8in1idro
bFQ/VmfMpYYrlou2PAunsPVaEIH85ih+HJQepBRVDfx8CMsctSV/Hog8KUIoGD5MrEsS+yGutv09
5q8eFTdM3Csmkaq/jzmuhwYK1SDBAroPvYvadkAPS3/e69nzp+Ga1FR9PZjcujxpOoIw+EMd77Zg
b84vXX8SffbLfTI4kvXd/PCE2VIjKvRJ6vtPwSYTzx2pyVjyBXbH2VwR0oi8WIA9VxSwxmK4Tzje
miFwK0Qu9LExILcBZsxU1Hq6T+myaB0YIf3hwYi7FvZE6okNsoazwXDlrBPnRDNOCC+rR7Je4InQ
Crl3QbLqXbjGf/zKV44zDnrk+Bsfg93YDrQwP6QdeffExBkdG+QGG4M/vBurvvPsetdbnz2inIhc
Ikn+x3C3lnxaV+F7nIRcpGiAqmmWVoZs2O3zVyy0B6+PgJ2YvQpgcTJptjdEdd4g4JMIi7yp5ljI
9RDv9Y0e7ptavGSOEpK2asIkVfGnoOWZCTVxbRgTRmOUIJunWFO6BHgUOU1RpDlLUP8D07+slZH3
O6Fft8XIZLJRvxxnrnELiQ//sN8Wl7mPVP5MAohCz8/Q1FR3+7up67jjRab4Dmi/C52lzwgcQNr3
GZVEJ662LpFJD1HTy1+4y/9qV1djU1bZCc74tAMtbc+Nl8SSKq0rClg2fwSTc+nV2Xo9LxCgSCsJ
VU+n41s+USYWR4LrjutU4MvGCdjRODenqnSJA4GLVnyBb8DeZpI90QzmcqHmUocfUIx5hw3DykMc
AFHfdZVUffpQrz5P/vEaSvWc5Z8Bzvzsh/JQQWPzFocpNPORteOkLfIeI6kjkbVeJGYJuw/ifqud
6cciiJ5x1FjTMyIOEan2gNk9a8tM91LSMAN3M3wFGpDzu+GDzsw2C3T1F5F5C5rrX5q1uOsQlXc6
AaUnG+7RsEVgxrXTY67ZnhoXyhzANeOOpPJuWq/PG5sy9u8L1BIqcA9jZcu/jP/Mq3bhJr+e6UR1
4mCtH18krclJailve7pYEyYK/qZ+X8Wq5YGecYlmbLfmhxxUpzSLzPysmqqxSvbnN4IiUjNKRXZW
9+UJpQPNGJjZIXZSK1gbRAZopbmU/DjLqmaBTSSjRlaEXIRFtRWPJyhGJ3N4eeFgRxltLoJ8k+tD
B1Pl/t+ZdsCeNCzgmw6eEoP6lGY5LSBmgINiVZWn1TkmC0fuCVIpCEZLXfsZwdP7Zz6iwRtPnc15
0BQBkogJ1kiBnq18EUovQdUPgzWpjp75Xdixi2ispYEJWl7L1B7zMOFrsrpB6vIhOkhfsC8ZcTxP
U+Jifz+2GiIw7GciUwTsyFmbeAx8pIlzWgizAgA3WjYC0K5cygD8lRAfJ8bJ9ywtnXi5KA18p2BZ
u6lhjKKreKfBNCUkRmzfwzog1B1xcG9kFl8noVexmMc/+n3PtKY9phmDHViU7HgSTAIFdUDv1/Hi
lami/lNeti+/F2sjPSLA5TR0XkNMaxq3gfnfw/WW10F0lKfX1rWxBp3I7MLv5ekuQ9FzL8Gw7WUa
BoKnAuT9jRRAOt+/CRQYhQnkcG0EAYBpAfXP216p1/JKxQitlWw7ruo0pfSAZnE0utFO8jXQxbjG
sc4/uCrz8oTADi8d09hABxFEWPv9ZAXfBHFJa4RmnI1bTR3j9w/pEosr0muoWDUJAIg1/6VkScn8
wiv3uK/mWgWlJ66UlOmtr1hm9UMlip5gJ/Gs8Xy85Zx3cwrXNhUE9vCZc5Q7TYiVikGiTXXNO7Ri
NwReDdQsN1oLUmCNVT5sh9PYLZNovL7pOsHQsEzPiVauiJWalEWiUM6PqcWjylMwZCHiCJf8VP7w
GXHfZUDoRlBwtVztLeVnktU+3XfJzn+RQNBMAOQQYmnm1auqFF9/S4Ij/zd/z3TbrzPZRMmBoTU5
q7183xuId26KVjkXYixVdRPyJqa+tEGh6npSeUBsjxqKFm73JnK62diIoKFBDIJl6Lli4rXaXIRt
ABE/ITSNT0a6VuGt8xABrRZvkzxxwnKFSLCYmd85p5HNbJ0uErkVs6gA3Vv6rMLEmaVPLEfylbv1
/7tXAXohXbYTKAzNqb7vjfat98fkpvbM2M7OdpNOBTQBepdPG6ukCAqRb70OKY/9qWkfkbFEUZsT
VOdBtoRKX6tJ6M7Ah/trgTy8f7MiMkmr5AdWmbjG0XvBIliW4dW4UQ3SA8pHZBAAjNC1Bep5QDSQ
wkY2EdFb8vBCVfCjfoVR3gc8JqF1OClazushIaxkKA9rYgAZgm3odNtnmWVXix7kn+F+BbZddvey
9a1JYxZ/I7OPDWYHNK7xRm1oEEb2JSNOcgzjbaWvtF9w5uUuJtos935tE2lCF+XucyR+5FIgeLa3
qfBvhRumF1nLR+ucc5M74VTl7KMDIRgcan5gEdoYO4fpEUv2eMYbaahBIAwoYVGX8fKSTKMkTJux
Us0OGNvA2bIXWtbnfWmHSqzB4cw3lnedW0/bn0wx5uT43ph/f2U/Q4r3LJ6pvCJa5PclhjxG4+Ka
VDIJy5Mhpjn0tTyphT6N6Ck8r3hdiorPstBA40a7dLbb+e7K7fdRIEBDRcU+K+/wUcg7US3V3N20
7qDQoIhTn5n7HrrVPJbNMnnuYgBTGZGhjibF+6oMH4egk8YHa7ALiSVXNw1qjXvjD6y45rdyAAOR
qIbyxdz0zuMEEr1w/0wA7qs2uousKOa+Hz3XOyjr+W9letK+rZ54zFnHoPMOSQeoFMlVqwOV/RPa
fN6ZipodVYlw8RVjXDPpbaYyJF4xRlUVYlU/V1Pd4+AQQk+wkT1OucLk27Zf7gYkK+u0O/JS0NBj
8i+wDtrdUdCmxDkYUSFqTQihli3buWeAhPhKnpy/437RU+ap+A6w9yKnc8+FU8JlzV0I66Xx2MO9
nRJQxbqsZEjG/Y7W9chcOpdAZL3CZeQRkRUihsrJC8r5BC34xeU9hH5hrXIqXnYEybiyNd7X2/gF
rnmw65uhhpNsyfBt1nLsxUtCDOc/PMwP/Qfdxm8gVpBvc2/Z8jkc7UaQF3KA2qDeEGE5LYbdNIM0
NJN0WNpgl+qtb7iO/81RwvD8gfj2VlGFZIxvTpGtiqLy/I5g/CoJ3aCJ66wH5gtvQ3Y1tZvK9a4S
wp33ccUP92rfGy0xnQDPArFSwxkDMNAHYUHJxdOdgS2ZjT/+o2xbl/DsHlejoTBh3+2pZclCXls8
qhv4hIr7FrVmn4BZ1X9mm+Be0+Hs2+VsolT24D/lYy/cvjZLp7rYUOjdbJgPBlhFRQwtFGdEm0rK
65Wz2nhOSBuXSi0sQcSBTWYd4v6boUVJOlxhq+8ldK1xcCMIJBkwChQmWX2AdHzMqcCrQwZjtf2c
mRF8PFFVtWG2wff2UBdaIqXESnjszn1+TZ3ATs8MBX0QPIzB0Fu8oBhE8+RZioXZUpnVxmD1GDV6
88h13WCwt8Q/RWS63Ffb2jhbBxE+/gMUtTDMUjNgd+9RlVBzTSCkJQ8mqDkvrMPo+pN/6O0+Gplw
tEv0ER0lZiDIVr299NlnqYj4xO2NlUtv1IIzlZMhHBEG75ZV3zK+a7e53nIekjHBJGvIn5KAAJHK
kP5ISaVtPZ6ILJfKWKcpF6kPTjQmyC6zw9Ntrm+6JSEmpDy47iVS7IgcfqZNdv1OWaVaINMwhuNZ
KKbaCs5AA+lbQ7D4+w5TbW2C+6ImBbgBflj7mkm0qEcJx1SOgy96L9PIybtTLby/WQa3FjtwqRWA
ZUKLIJ3C9LfZgy6dDsf7EgDO0hLD+vgh77Ip5OC1cJk+1J/x0mz8PpTgntL1AHHFzGZEYqKwuZXK
B2AScikIdue4Q/HxxUKBUJkERnyYklR2edtjkWMFik2+LVUzjh2u0jaUVtAuN88RZeNH4kieFm2O
XMi6UPE6Uq0eeJb9MVyH1wIO7u3i9h2+90k2yyEyoxGboMpe/xOLUar//sY/tY55qDBwDIU1PEO+
ao+O5F5M/EcIZBHgv+M93fzLWwf5k3J1jhLxSxhvasRSAlbZyRbiE+AWrhAhSqzr5+nFELsQjNzO
3/8nJYrgSOb63Ud/xMXI7LetxWr5q9sOM41QSuk63I9FMmW4GMdJg7MxCCMRoVyON79wbgF8yTx/
iMtqqtPwkH/zjIA+/wnDSWFDOWJxeVakOn3w4KAu6CyYod6CLfkjd+2ZKMVCfBAK7bCybqYA9Zv7
gPQj5xvX45zjMNlZ1ktR+x3gTaWgZkns4WlqaKEwgESoWp9UDKFiU7eVoP1UGX6m6GkY+fP10X9W
uRQFEo2njxg9ddUYaEN5v5kbLhxqW6jrDkx2dLqIGzlUzspnJfhQgVo7YdRMXm+Ly/0BGKPdyXHd
ApsTyH+hoWbDl4I+t5eMMO/VGqp4wTgppaTdLdcFmi9v6CEPx06P9gF6B4GUf6RJfElEvAR3lFo2
NucpHouyBySN9ZPd9MuSwsTrx7RyoZ5kkcmflW0fXPVCfp2X2IVKWv3VZQxLP/qMdIA325VYCIP2
EP+2g/2wnvT3qYWSxDwZ85/blZ+86jlsLJFq442y2JU0art5cNLdyW/phIVloeBoPfUEcR9uDL2Q
atManax5TfKAktcLOE/HOdT/Ytu9PnG0S2z5LWkCaVaOfMCnPSocxzNNyUvsBG1XEMA55vgHK3by
DAEOhX/vOXSReV7Xny9UWOYu3ttrgGvk6WFbkQzNqvmx1yIqWBDWdXEMKtbLy1sqy19iMgPkC+YO
RU+CHu80cvrEpBBWgmQxngrwLaxcheGFnCLZxYFMRIU5LouhIQZ3o4BH30nrBMX2pImdMfDMZx7g
AcSe+RCs+N/xr1DfYRAk5CsIqfitU7m1a2FYe0NaJSl1+2FRGqaU7lFRZBXfwe89D0REYzMhApnS
sYwRBLzXBjDi7+HV+lxv2RgbLeHUwelG9uIV+tAQbaR5JeDLndWLLXEFRMXWluaK2JlyeMhUtbUc
wkuTDwjQtR+1jTQuMlgrVYq6UcMyiFjk4h22FbAw8U2amGgpoD58GTpZeFdexkZhQA7+8gPPvCG2
XE4MzU31GNHC9jsZenZdYJRfHaoWDSPOIwnCq3N+kKiLy0GuJIiw7htnarzvdVZG3d/EpIs+4d7W
3d5gwm5ubtgC8/SsFkp+Z3n3bsz0j0l09cw/jSNfTU+wiv1SNTH9VOASt+wxiYUU2dFpfVU20JFj
tM2airH4XpVnfdG3Y+uz+mU2mpcae0a2/suWfsX143X/5A9Xgo3KwTYE3VvMMjnPfwb2KFwmopQ8
C7Cl9s83a3ST+BZYj2xZu13j7ZAYxSQd2XUC5wdOwswVgNV0qUK27ZW3LNPLL4hOXrTCu7kUJEKa
ompx+UluQ4+3zd1ZQFDG+nP8UD+IWggSMZkof/eFSdOAjWTl3JNYYDSjQrEbvce/QKTn2Zzc+hQm
Iv2qaPwaIupIyuOGIHa9x2aFd8hWeD7ZYW5OXQriUOucl7pf0TI+B54QjEOlgNaLxajoPnXe2llf
gH7URO45R/V1bLXP9Vh6YCfdiafHOUncoeqtrfEGJs535ynklFjlEJ8coIVV2l6e9/d1hORUNBZj
wDnt+n7esWlguy1JLk2iU3d6rL12w41b6BNSAA4RnB0OTH/fE2To8imiGQe2BdzU+8xpgRN7r/26
xyLXSIUNAI77vzoL4O0TGwl3LBZ3mACyivAhy+l9IC/gMZSLERTowzxLPhVNm0ESHwbq91TJDm5X
tEG4gZkT4L/HINAjli/qsyVt4/Xjc6glApDPTNz6CFd8PyGIkCroVwrWbOU/5EHCrdMbEIXIII1Z
+sUCTuoZqo36gn76BL7YTWfAYbIiuw+gALg5FCpSO1xaTuiflRYS3r9D2aBT+SE0Au+Nl7bVk7kq
6HyOhu7ruC46HEtsv3KgXM2lp5VnghsVXQ4SL2XavluB4Pkipaq1imlY1fj87fVBnwoTloZNuFjK
OEBnA1Hcnu42CFt5TVojGtR+4ZtJq3bxSOJNJBgzdlN2Q68elAHpv5Khleqa1tySHd1ojydsUeZP
DS5n3wiQatQxMiMLp2wWodrXCyG66Px4eFvGsbSEPSVPpj2YC+GgcLiq+S69z3H5vPWi6axgKq5T
eZannA0N1ErqhHpv1UOEr++7STmXK3EkUSZfJ0wf01ZlDow6Um0hHrCOw/F8FLIJ0exNLWSm8L70
+LMqvAlVz/ciSiIhLQBO14jaodkJsHjU+F5o42TNnR/RK4VxLdSAxSYhNDo0wgExtU9eQQvlkma1
C5gAx0HIQyI3kQG8NbnKuStCHE94624PazdzRGfKfS2WkcTnYUDBNkauHj6cJBlTSnw7sj7EPWQg
SvLPYZgKDp/RlIarQTiFoVWnEjMPUhIyrHo1Z5NrIPHJ/mrZuZ/l7pyBakuob02mnZT7VlURhCMp
n9MnytLaqP4PubMKmRbCmHmBaOLfOQOjtJEVIMyXJLCKBIDKgsz9bXD7Poez4vqOKdYh39gYtc+Q
aanvkyjkgbnLqfC+tXMQdwnJiXjPXyCfIW03We2vLEpKKTOOkVf+oJHtevTtEEG0koSXfEfqCmQa
+1bg02wbJG9ZxLLQp0P+Sv6mfhPOCwBlKMhOMZfVumgtltgt3oyj756H7PUWTXYEbPpeOlrqZwDi
clgFZpR92MkIvYR0KfD0dypEz/+QvrzoKKVdND9lUlW7GEJNlcDvTUAR34fPF92vx72tCQSJ30f3
wQbR3bC2SWFueZLXVJJ75YfViWosXu62b76lJQFa4KzQCAQoxr/N4CGFsPTYmfifYSnuoH4VXSO/
nlBu7yaLJF+9BhrCJUbko++/syEGViJ1LHLTdCVXvfLxIomNS7sWvg5Pd05cviQhYdNHc7kog/rW
eD8KETbSNWQmiOfgX9bN+IhCVTSpHCEz4etn/cTDF8yH70rNsKsjTm6yqqVdMy9TxochICCUmd2c
hQLHp9RQMhTOXeRz6+9Vi8gNVts0Ym3jedZ1KymtAmrtYjTEr2Ftdl4xTkbBp53DSb1XMNFA7iCe
x0m796CjWPgQgM1+pOs32FYa+bt6iHm1xHyRhNgp+mRDyuAKhWY8qpM2dtLePiADSzzoziiBWvUl
fAf+SWayysCO0VBN+NQIln1kg+Vg6d37uK0r+umkzB1YMzbsqxjJWiiQUGjBkV5zP+wlpSydnUBn
Z5g0pBdd1jtnmx4v0g1E5ELMgSHaHv39gyTfeAqug3BJDXXMicjZ8NBwWQPsHka3FJhxjawi9ir9
pm74f5+Hq7HCkirFdEA/PGxb6yEz0lfI+iE3OKclVK/xWqm7Vi1LFZPDzfGRrFHTQNKozgSbPbBF
5fFlLPEt8VsVhAgCrGhJBd7fIliXrUjq2NM/10Ccs+X8wuhY1cGJRom3ERY+pPqoyreQ6BuSMW6d
7zyc7a0w7P/9Wqdtfe9O6te+fN8GyUsH/DMr1/ZHTDM9f91cSytVB3TG9OzAKEDWy8lUSd/Qp5Fo
UXOn0tQdkuUBIIOY7cEayFUHJN2+gpyVz5ZZY+7CGWYuJ3Viq6bHMdpw86UC3WKGHBc1nBTriaKc
uiv507QJ03/hFkvPmfhszKBJk7cZ5pcZ59Zt9BSxtc4LSxuoAlRu8ulEy+xW+2zn/9ixc25Uo4dO
Nz+KsxjFBsA3AdIQODJP43mZk1sujHmwxM5lphnFB2SNcKvvZxHhiupLhoQ15giO6w9SOjD8MQ4f
XOiyp7/HR8ilAeLjaKeEznc9qt++EP8Uw6pSA7Xv6+TcBgqUirGztfjU867p3kjNGW0Xsrw85bes
LQPIvhIGbz2jiXW9kcrNWJdbvoqXGR2Nry78eb3k61vIHv82JX3mJC2Ygrck7hrXbmQbY1LYNICe
+KMxCCZQaLC6OZZ7nY4+zwXv7MOVdedGonp5rS6iHQ2GTOyXbmnW9bnbcB99Uk15O+NdLp/FbPz2
Fg/VpbolPToa4Kq+tOKqDZ6+kXoxPYTGb8Bge8x2GL5cjcsBv+YRvWxns6fuu01JEDdEAJeJjHPa
5lmzTKwyOr7aqQYaDsLnJVmTodLoHNCiRkC50qMjrCaitZ7XxoXE8EF8Gt19tCGYH9wL5UEMDFcd
NeMhinfLmOM6iE3JrICq4mvD9W/CrbMlrehkBKCM6KSyIGCzUt27t2vOUM+IkkKVIdzK9x/qoeU3
56Z8dyM41aaSrR4l6FOUmG4rZbzwcXPHrmIS3zxy3C2VI+KEx9EHqsC+tQPH5/BPZq+2ZpmgzTn1
Oc4A080k1Ic+GD9bJ2eLIL7QV3N42ljSqnjAVNDXWBFkScMKTsn2cM5cbFnykThzQIJnuoGYdyTA
6Y/5/0I+QqmCsgAhjYAjQspeY8NYNYwe82Djhn+BmUyOUT5Fno4MQR5sXyzcdtOSfbtWyBBXnOlB
Yt1PsNIrYmQbvx7GsOL+pfj4ICFFi7PxdqnLY9iGq825isy+r2AxkhXSZm4hG7JHvWRjIG9HqJhK
kxIBc1YDYHMMgO1Pecs5k51x0K3SFm1zxrGWSFmgIz70RtO294b5oNybUDB1c7gKhq+eDkDbNst+
Vpx7Zt/2XqyW4yWCSRXpr4cjjYKpY88zI662Id5IDqFFJm7zURapnHL4U1ztnwMoRtBtj6dAB26v
FvfGl425Seu47LO9Hnx+AVr+SSbPoZBs6jNnq6vsP/Wcbkwqz0entNXFktB7f6DWIL1hI/FX8hH0
uP401oYNJSQBwjyB9nUql/TI++LdmN30r3ELwu6SrD9nGIS1KAwu2wXdVx8YHMzYJoA4ziSxHqFZ
3HjVmRMfjUzLMKQbjWydrasjmHMOeuY7gL4NSrVtDgShbvPbP1OaIBXVM0GhDVNEgO0CYuv+WCgz
83ctZYGHJ1EBmCP7ZGPEEjKN3Pn+6kXS3NDYzyuMqnlAE32K3kAL5i28jNS7/LXvdMzAEIBXGRXz
zf6rI9DmonTXmUFsaC5XuYgPajNERfRxCfY1dBU2ks01EaGnXR9s3GzwUMPoCakbSWbWs1CjNyk2
5Ku95uBapgDS9jG3xuarM/RLexwKFnXheyCw0gNZX34X3GK2nG+A3G9ESmxeWWh78yXwZYm7lWzM
duOPlAU7tdxIcir1RsxCLz+ZcOEWEd1crxhZp4rzXPmGP7lceL/mHeyYF81oVplUh06nzX7NW3rj
LiO3jmuKvF/ad7axWCvP0KopdQb1sagJpDwUyNSFNLzxxYgzmYsj6MrxMpSSOlOe87HYuT4cwYay
r46LYmzsAh1Dy3Sz4dBbkVsmMsZVrvPlQ22CV8Dl853JgtXtHCSn3YF68D79V+YxozgSshnNP+8h
rB6i4zfvTT2FE3YIT6nXjC3NHJYLc1EuVvdR3YubC4bnwii++r7d7A5mggPm6TApKl5V5e3jgfOb
y6QO2546ElzudpOo/AqFaWrg4YK7YXpTnpq0YLIIP6m17h2xljxy8sSGJ1jZXuKNgTuXbyZRzkK8
/DrPCg34YqWbQxD/TAnKatZ4vzavW6CexgAo+TqPGI54j/8YMdW5tQOrN+b+NHr0OA5qmhcfqhMG
PrFmdx0v9+ulceLbw8iM9kwf3vEv0fpAeLQbjY9q+MuIEwd9XUacZD5yWXpDg1S3nrU3qFd6T0on
HMk5jd4gzVTBh1cwL8IqmPd1iCAkq2FieZL7XOlFyHyc+qAaL7pS6VcaEgJRbwWsL0qMz39xWd69
Lrk4c2w7HGezTxI6W7d5DbHuI7Ss09PD1jNqR3mF+NB7VFydfgo3W8mh+piJxYzlYgL/nr6Uv5lV
a58mlGNmJArpUOFwHjzIgUCjhnV5aGid+Kwq5Z3av1zD3tV3qnppd3RHAHVkiwpiwn8ihmPNNWh3
SmQ34Rh1Be0FHlN9ZbAmQK5j5/zuWPxCmhbjsVif5a71iE+OMzNNZQCWHWK3yNdLfF/S+Bcvor0O
tFGxVnDNFUFZ/UHEpgVs+JND/ZhKAJgz/gXFS+IUid2GuBgNifL0oYVxXO7CKmR0s40ArAuNv+2J
VUa9+9qOsO0J7dsMVT02uvZcFnDaENv/a7zh34xq24DdfAh5dpJAQnegWxlIgYd4N4QxX368hWMK
ab7Sq+jEH5yErs43oueSM2tEdhq7UR4AdYAEkV1iyo9icxzKETkXn4qiUE3m2lxzo9o5iT/yVSey
qJySOcxRC5XBTWkyRUnHghNir0BPTY6HiRz/1+LlPgEMe/K/VuRk69ovo73LsF4v7877E9q5mdM/
Djn8bL+nesYQYZXxQTxiFxU4bcBCO2QRuOXdW7YaFn/NFvpnouZ72CWLjgTKsEcoY6Qz98yTJwlg
jXw6SErexMeFIt7KtB64JyJJFpT2DRSAEA4jK30xrLCLVEA0RtMgNgTEdzS0a9RmG+UkGZ0arKJ3
YOZM1aJCt7pyZ6D0NRGyq2sOHaoosDz2oQUYw+5clv1h8T50UEdF1Yb7iizpUNq3hcgdKKZoahvR
8dMF5aYnIlnZXjkv4FLMnEbE2P/dD2wNbCdvjrD4xXXhqZdarCxLPS6bUJ0iw6QNcHElmuz5PUaU
2F1+WOl1EYARgU9DOz50wdvwb4ic6dp2QZ9hURJXzNh9Fn5hZ1LTxztg92zXx+ngNsa+lcLWE7bT
JDwhUptzi/VorBdmluQUtLpP3xQKcKzhlf7GEy8gR4/3e5iDmNjtdf9Kg+tlocUbsuSY9SmbySDq
Zb6Kf2zaGeisDr5hl58pz6EJMTCjS1tY39BIInXcrqRWnCpDK5H23IQ18EmTuBlBrOAp3dg1F5U5
AOayzNSVAT4TTWLBB5BKESf3JqgNFiCLCifAJJMp3XDgZwKE+J8lUj8BXkbeRIagvfeWm3MUmktP
aFEhewE4K3DMdckzyfMhDnuH9RovL/AUNYo/DiPb9m08KFfXXrF0O/PSAl4Uzut+7CXqCSITIe9w
dU1SlJXSuXI/+AaOD7pIT1Y2faak4FOxBaIitSbRuOcLRmWAPNylJxWHdpR783NtDxEdeWRaHslj
CXv48mgxO/eh0bU4Y5qBVh/p5DAfSdJzoxa+IoC8jFExGi+W1deN/N41UG/1sM6pfyT+Lch01+1Y
2IxYayxuRJNUYDgb/OvRuaxpXpsUAFY+mAg0VR1IIEGquh+pL8mxAyNiAP3C6khNrJwhoyU6jZXp
UsTgprdLCoUAAVZ0xRmtcT+UH88rj5MzsFqR2A4CQmGbxAYMBBl3dBVikEVFlik69IDa0T2sfUOJ
wQmh8zkHPns/zhoSKRo/17QryW3Bt30kkiL9RZKRBrk1DPdZdn34fYWSBR1oi/Ud9yFycDks7UsE
6BWnZZVzlrhxbSjyd7o5zMl0OlYTdpBtsywMV/j+wiH/iqCUWWO19vwLYRyrRy7qHBISYBwTTKGH
QbDGUggh77t8GJ+iUjuVcY9ZfZ/kFgXg9XbqtMqkiYSiik5CEbk3rh1qZjKzeyY4FGcn+fiZ+UBq
cIJ3rZE4aCfy2wmfQnCE/845TYh0oRI64Bd9zaqJDzlVwfAcuvM8Xn0rPdRaAETFuL0ZKzdKuDtn
5Ls8BhnL09H1GkSNDhIubITeiqDTXAQCtqWuaaLhL1HgGx103ol6Oy2F5AH0oZZqIO0FGLAWcWi3
Z3/CnfZC+9bfymsnPQdcSnot25i8Bwcjwt4HnyiiAyx/PR6E3o1SO4WlMrclJxw19PgiIrNoteWv
QHGTQrICEnc7hOldaBbeE8BrmbtEuCvzZnhnd3gV957IkDAjRWzWtP4psIFXsnJ61hwauWyFn+jY
cZsI7U3V6dgzVH6UlLIBliz3G4nMoRYIN2heTUiVjKPfRUn8rexBF97HMizVVo+bOFfwCmOevRcK
wHj3R9mjLJqgBLyloIeZ6aNT/R+bdYVTldQyrjfS6uZ3GMItKKSloxoQ2J+MAsZfvStx35tcgPds
JaKr0A4A//Qv/hhZQNAZWMVkG6+OTClEWkWzyAzCeh26tsA/RV7KBT6b4z7axh5WaBrxdXvcaqGM
x4hLbyHWQWgCKKAx66+QX7T90fOdkk0RVvl5B62xsoZ0ox2dJJ+UOWtqicMe5W58S6IOyx9ZnnuS
mVRu777a8aU5mdV987H3xnYlug9UXSEcSCznTkVxdpZVId2wuK4SPLk/rEumqUusTHj/RuQs2y42
4VfZ91MUNoc/jMygwZgt3/L1I/Fb2tChTuL5RXaC1tsEUb4ZXa8f8AgQciaLKH+ZnPktQhNtufrj
ID4zvy9hkPF5fBXvidcTaXa2xGk1K7Qwb8bggJufk7geouuItgN+cogvsLKkxr/51GUvK/0xMcjU
4rnwBLVPI9MVx2K7xHjizfxiQ4EmIlBCyjAOBztiqxvnbmJUOvj1DDSMjwGsk4ugZ6zEXW06z663
AlH5KLVPo5CvfvyDhp9PfwKIzi3jK7lvgKVPXCfOz+2VmgjnZlcDQlpxf5sOSytfY0YCfMBOxdec
yEiCWGLjfz/itthIGxqpdTSN924pXaAEk8BNSojxHckozuT89zE6+yCx3KCDCuKVw90Lx0kSXgq1
jRBSCG8l/hsD8qQFRsW7YrWfP5eO494pmjbpx2+0zxtGtwy0Bvx7VqcpzchwxWOyI7JTfaObJPVU
XLQGYzttyPox/v/9QhtAW4BYgkf+Q+q7Et4JjT4lBYOwG65VyZjtx7JmyTRvQ8nPKehKv+lf041c
ShU+e1CfjuntFnfcqwfP1/ZxC6UoFgAB4wEXp0FwJQvkO2jNTLLPpnZmKv5mLxTa5z23j9lVGjWT
RkYWebZgtUnEpLGUaJ6x1nZdd5uNL6EY/9iXiNYcmHRinLU3R/3Z69/l2RTDc8teanOccogfZtaK
rsx2sl2NMlHmkyLWWV+QFBB1B7uWcciOZreNjZsa967BxR21kjfuyFwEIeBvgRe41b1sNzz8bJNf
86KgrZ2L8VaEZzOViShE0tBet07/ypAG88kaUolOkfwQVQSJo9TOZyfuC0Mg6L/VnQSsSPs6WBS6
gN0ewBy9k7ruQsxXAgSfESsu/q+YEjHyQTHrQEVdwC5xgiFPZlv6Yx1qQqyrvJVbIuergfa2PCpN
MSCvAj/m0qmdt04Lpc6szFa7SKJ4gRLqCWJa0hL/JE8aHELw6CeiHouKWH73Q/DMGY08OAnlWeGF
eI5hYKiUTGlbygwgky1Ocuw6j8NLXkJtZdU9utiMbZThAdQLk4RuFU321v9aIFAaPloLnk79ZU1e
VPsFLo5KdajRnaatwtgghshgGPSARihpqSYv+zvBE7a7q1Ih5PwYDkJzGpRk6UZ1tJXcWJ52aRFw
Qd1VNbaM2Ia5mc1NFaVwjAY2TK8l5ZtbbKIKCSDLofvUd4uGs92eNejNJ5LbWWRa2XKNjWG+V9vA
2hviewlMQbibg1qD/RJKyNLzMfcnh4Ug6UoM3OCwA5w9t6cfebTtCxeGJHiPxkvKfny4Wz5sa2Vs
VH02xj9k+dQyuqL2hT1LelGdEAfd0ZTApkCZBn+NLSjTfaOhUFH/1IqdIF5YC3dKKcpFqMmK7R5j
+XOsWb5EiV4th7hkI74rpQrvqYhfie4OvU5Ks0LlzJwF489ZDDyjUTbhMTaSsKoaEuxIuNhrPK92
uD9V2w8TKs2BeMM/wBFUPswVoZN404/rvA08dPDkt6bkb+CUiNl7BF6gxXD2Mj/bSDwouTb60bBv
12CtG140Pp33uJZkF8AwaEuWZ8aqU/F4bBadiWkAKIYq70uq7JYXGth1vwSSyFHX01k+tFfIunGU
EJ67oo1gfpWagN2OPebXdFHuDz7u15HuR+sXx7QZd0rNOplbHvxRCstIdk6SfM4BYKC10Ia0xRNP
JeA2QaUH5wvOaI3zYyhadSlk3sROO/IxJthQwnCaugdvvaY1HTCQUsWKnQ3/p8PIthblAteo0Cu9
a7yJ0oLuMJZxcC5FVH9pjP0qSkANuzhMfnsZ2FDa9auJM8NjJjFg+6l9VToqncmv4Y1T3XdWSzIv
5cQ6fW+0JQlKBa30ln69FcQwY1H50Dzw7q0ZsXAmse0bGtkopP/ZnGnwxfanbdOwaEtyVq+xeOAi
/ETZzjBtdf2BJcwovvakoQl1Zf4hDz4G8Fr2hcP8QXZ0lEfoVgCwEhnWb8lfI6w9/2R0TG8Qi8XR
Lh8aAYmibxyzhaR8rOKczsiEUWsw4/waIIvw5LVjOf+ONrWJ4vcgJSqGFKXxZSJMmpPLSqqQdUHy
6+wdzLtHG7qlZBOonLAHtegO4ZKuqwmn5O5BaH3CHFaBuWB6g+ZGCmAAwAu+UHv8SmXcKX8ybTBU
fE2PtQ6rOFh903rWRmYu8xDsXtwAUQjizQtf1QkiLBALsxiC6wwt1ncfxcAw8T5gMPkoHm9XNJ7u
zPp1DfRvgMAgp8ybhz8Ii6Ik+K6NhFuS+qyD3/nbpImfPSjJRnXU/+cHQWm6JmbAEdEfWV7mCSDw
I8YLrBc0/UNAKO4Rvgz5XGc1ADOOyxeZe5lqifcf4yKAHNaWIeHiyQy6+mYbMIhtZOQZ+V3mmoEW
0JaN+7k0wSCFg8v5+ieon4kzOTpuIzPQXESQDK02TXQIkaRYUTsbVuIlE31v+z6gwoU5Fh9QwTrW
PLdJWTWRW6UITnoT4fu6oLI9w5xCKpRsdBc0w+Is4NvclpAepwAsEwoknkqJZGhIG33nPDMnNYo3
EXBDDmxagdI5oaKyy/OBXiL8p4QFGt8etkjBDFkTep4cs/Iq6nkBcCX8/BQXEO5xK8Pr0+lJ2BPW
O1PQmGAdZbYlxbt/7vKXyl6LPeborhxiILrLhtkOi7UcwBzn59BXBx/neRbm6jyBVcpcLkzwAtKf
IIu7WWiBQ/DxK1Fl2n4XueQV8icSqussr8kOMOUpYMwWRtWc+nF59iHGZSGIvj4+4Eoamri8GNSu
/xWZlUw0jEmRIHnB8UxPdVp6deK23eLz80LJ8jUeFnjVsJPF9Lw/8Tw0B9S3Caq1Ht2PnvOWrIsl
7fgO1ZOO2v+wk+ixwfXliqQ1dKC8TYA6ForVCyb2hcHqOYTXaluGaJodr2ebVcB0FYf1xzNNr6xu
KDNTVhVWzvFKfTCN5uSgkfmTCEaQCzseRySFgwKW/hPcq4ReZtSKpM7Y749eynD9oO+V4VJSfEiQ
VYF6zNTIvbN6/P1VL687XW4TDmm4fiPT5DRxV853OFrcr9Y98PyZomKN2pJlxQs/hCwIkavCuXYE
0xAnSgSzaTUMx0+Sh608vDB+5y1Pz+Xgvq+9headzS8NCKVlh1h1xIEilT+5iFuYOHBgRobEhdXd
JogauOnYrzaNzzmZavU1V8Z+C0tst2PnPTDFphVKoJ4nKd7RRCMst8Sj0WSkyqwbrUaA310X/Jup
Qp0xYjRdZlD6DaXXbvhUUf/b0uyY9WEARddo6oFPswghjRt2gvNJqBfhjoMtezVXq1oMK+oFExKx
v7tDZJALHWl6FRbSd/2FrpcnUabZTf9f1GXMy9KxRpWsefy5uknC0zIDW8Vc4kLTVx1f5pImmFCh
yAU/6uPkMkSAow8ZrEPc8wgcjPmopXtjnYFwBJM9Xv06ONOI2dDmDcllWkrcdeIt8606Ld0xc0mk
baVNVWs//67Wb0l2PKOGvvglwoISzE6UyMN8J2YBxZK+i43AaA8VZrb5OwX4/f9aq6QR/nVpqji7
tXByZCZ1Fpnb69h2woEGPXhDSYg0KNDbdrCKu5c+aCeQP3BivPnyCN6p1zktGKKuuZu/4F+gQpAV
ezjwgOfdzMUzKpCvx6rKjsefUNLV4Ipqxtenl3oRBwralLFkQQj0qwLdQdDwxArzQM0tJB90WqUP
fZmc77qa6JXJCeaja4Ij96/rRsxVk4PgYHjQA1hAPE5ARoDSIR6t0mKZ0xQC4ZEKsz2rx9/DajhV
bThqTS7ouhVC25/nsvoLZeyDodWH3Fthc56cPzXNutkRFPlaMFuaZpik3MtgHDENlR4azU2F3v92
CKcyJyHmfrOak9jA876UBa/CprBWr/wfh0gh4T+L+bVsJ1MGlS2iZovHr52zwWPAztyXAZ1ItJ3j
9oYJ54TjEX2zw+CbI7M+fSJO2kUgveRbun+OdtjsCBamY3j6w2ez7P1rv2/owi1fe3fr/gm56UVW
ERH0rKyp7BnEJIoG3pDlm8kINSU+7KIv0y/np08u1nTcD6a8UodI+6NP9NA/0I2O7tOL/0AKJA8t
kEECtZECC+Mh1W4o98DJhcYcRhAKRNqbRwv0RUdACPXmw4kX1cmNxVS5C3hjBEYQdZqCvxXNO4NE
NKi0Qayaw0yTdnlDN2Js2bZ7r94lYKgx+3KCOgxkch7tpHEMI4QOTR3K2uVJb3apsvDxhuDHg0a3
CnfWnRATRYIkWyevX8odzMokEVigbWHo3/EQEQD/bnFI31FRnrixpExJoTnpMDLTLYEJjQURr4PA
0CtdrO3JPevZpaHMGzfssxN+KoFAS4xsbNwirxF/rVruXs1EJp6TMbjoCcLZuNp4MZrh7sEPQM0a
h2gRX9/tiBmMMLw4NQ2SoRE+q9DEEzWwFxOZtmHMWRNTwLg260YMHVoFska5qMh0AQlD77LCT5qA
46jJrIJY23ui+wEg498ojt69C5CLcGpzNHPV0gkkjSoie2x7ZHGTtv7scb3Fyj15aN9vJUqcqvpl
F1UC4BAG5HPdS9xHt/rNXqIHnGW7XYZXKf/mQ9ut+RmzvNSqpPXZWJH2jQ5rIGo1MVPwr/WNp3S3
WRsB3ZVmXaPwhopOGRU/VDbzM+Waw+Bgb4HG5LkldWG+LJPuT+mkqfvhuwczCq0t2ns0TdYortQO
fDLbmnLeTJbCkwbJD3aRFp2oM4dhO9kqgAVGmh6VG0dBmCBMyftvTum6+VhOHNDD1E137BAZyrYn
A+jwkjsu48osk1CJm7h6JtkfzZHJ23ZwGFH42Md523MtG3oacGil0/SOFTCBYyKVDf0tvMrokGAW
Mrhz6YgVIvnxA+XI1/g2dAFW+jQZF2NTR1gKEsT7c3qKl/xUWDlYkF09ZdL8qq5lFgo4gXK1EpRo
39Tpm3IE3eUhnxC6cVlz4Wpu90QksO4fC59uDgTvHPvf7OVflHKCXulDs92wZ0RtQlR54GmJ4agp
PRuia0UmqCoaxXHqW28IRFxiKWe5FlGdxamlEstFLn/6zHEhcUj1nx0cHKNWWDX//AyviY3VuDJR
sOaLAuTdv53p/8zK8Hi4a0MdrheRl8m+72YPZXrHJyRVUTfZJYjpx1KXM9Ryk5oKuZJe7POnDZtx
KqVWdgQEYOUw4YE3FPwKcJxToQ41i3GWC7lvDhBu4lRO8Dtq8m6/X61RXY/YV7oZDXSrKARjnds/
iBwmUhQsShZEeyVWN2f7yG2y2vWCU3bP/YahRCl7porurtIEyiPFQdHGlhuQVqeyFyFb2HEC6H10
MHeVBkHQFTkx3wnt5Bu+TVEIXGwydZtimKiYyo0URM2GEo4niudvrTr8AH+9LXvcCR8cRRuxUai4
ucdVpn7MRhs0q4nwX8TJqNhLv4xZaHuYYKQcF65oE5s3UQB9ejbbaLb24HseIOjWgIdQWOKeTNdo
zqMey8OxGanzA48SZXCWkOevvWQXlWQ+dHDkd0F1KMCtH08iUgmi+4OZVHzQa+KvF9PW/+lleuYk
dXXZn11F5aSLEZ5hDYCL49paGOhDS3oN5nOt6URr20EipfRh2jte/WsYdaU0VxXqLmOwA9HJHagd
zvn9/uGXCePSVX5q7jMjWtuKB7FHNLQ0/t7YfriQP/zKx+EvOi36uX2GhbINkVVEZF8U9CV+Oil3
5oR2dKoSng5g0Htzi0oWqcVcOODa3y5Vx0MR1Uval/v8kbzk/5lqdOLv0uYUCCFzygn7h1VBb5Ir
3Mdoocr/jXthKdfj4GniyY71fsvNoLWUpKCxMhiyqscybmAezHQzjKwsi4epwmV7+NkNcsMXG1fR
KhO2hQGeE33UYRi7mdeFPqY5TZ6ynx7DCE3nQJIQLoMa4DzbvujEvQOA4hgUlJIGn44ct0HSYO4r
TRxjCVGJhmRnhQkzBfznQOc3p8XCU4h9+1PO4q/D7jzQkOHXzO2aEJUWfPfN4haL7m0DlKyYauZe
hFiDsxJkvUmUcJnrS4yVyluf8Nc/oYyX1YLMgFyQ5gqg5d6RlLuMoh5J6xyBJ5jS0grrwYGNunzE
1YM5mz6Li902IYwWFpq2adqCMLLf83NZ7GABJG9GEfKLJHk1GT0E7wm0Q7GNRzOVzx0JKA1Sutfr
uvTp2L/QnJyvUzbwQXAyuIBog7HW4niTAPbe4aW+NRYgBLl7zoS8diwQ8JVrjfdmfcMv8SnbxkPQ
jAIviTejsV8y28JL05SI+pNJTxYxhRD8H73uKqXcRW/QFMCPYqzNPP21KkzFch+9NceMRgm0WCnr
YfSXFhNZoXaQmEa5VKlK/ctRdkCPuMmZD9Ji6pxYGYPYZQaLJ+qjoiaqJrgLWoTeWAOpSgn4V+JX
H7WgKBqc9Ik9RjeEO284cH0vtknvQ3PaLvEBdqwGDHTPvk5CRq+4qoDRAJ7kjs8DQGKJ5mdN2c1S
RHL0FEmqNUiBj8//qi8Nkh6BNGKAN+VYEYLn/n3ZUUTDtMWpbXF2IQG3ZidMeNRQmyqS1QHzBeQZ
6UI9K7QvV9U+xmlZduYuzYf9tgVGVVt0Rs2ACyPV3bJ3/bHwg/uuY+xxN2ffyTzbMTM04jgdN8Uz
jwuNffm1EDtTnfFmEG6LN2Kt3bzIH8uVz7JrPgTr3uF4xpa2VYTpGf0kzohwGhp8MA/p5Vy8jNVv
jbDB4SASRPcv4Jbg9gju00seUNl5BcjSorkoolkh3zUuTZQqrNOlrQz2p+yhYVdWXv0cqykssbFw
9BM4tgl1irUi5mhtBd+DhorANE0VkD5GXG6/OnhpbBn3ikkhBazrdqZKXO+K0bOgUKM7Nz1LvzAP
UzFNstm2hW+BXBoRLCQ++0e083+NtXDx0M88p1wEuI8PJz5+htMpvzYlLac/xUu3yetIODBwi6g/
SZpK0eKWFbFW6jqPVrv+R3w598wUhtIpnKrhgc5UcVNzV1WU8BDpQakbWIHLg0NycqYAidTnS8yy
UJ17I1rrHtz3akq8y2ywYpz3aLPmojBDn8G+QqpF7Cw+IN2+sQuhrtUdvOBMg/tp0awX26E9wRiA
ouFUiOH6sQx0Xo8FH2fu3sBbxMxi+TMggW8waC/uEEBVtOKCDtL4ConVEXB9qgHDyzjDQuuHW1lu
sNN3+oi8QFjPB+wdyzofykulfyjMfQWOaB6tzcejbqtPSCF/XaS/FREwSObEiaki4tiFy7K6aYeC
qjvLQ8dGy7tGyXmMELHOCBKtHZVNPIaeqPnKAmaPSPfTsyqPWjLZYb5b3K53f0tWWwUWYEgRXMki
ncuWyYHd464CwlmS7vRg5xXiKwYPa5gA6kfC2/r++9jN6nDY/CjToYYta018Tc0W3gz+ShawYamE
YgSXoajUTJFvz2WZD0ESxSIU2zkWQMC/TfRwmW9XnFDk+og25Id4okZ2ECMMXurGegN0g2Bk9r8G
k6Y3HMaOtLuJnARfiutUbwB0kLB3XuVZzv8jNZ2XnRcQlYApL9j9UAEoMN0z8PMOD/hqiGsngWoy
sOE0lsBOSO3dZ7PO/g9fmyI83OqxsDziYeegYL2044wkWQKAfS86aYXtSuFsGMRnoLiHBQlZoT+k
/X8IXdjbUIvgo4ZnwnIkOp7x+M1TeODX0wC0dJECECKbD/VXfuIvWlBorx2eq8Wx9mgniRswevPG
k2eQ7auAwXzdGYawwbO6zLZyyY+lpYIKac7juWsdi+2p/2SyHeH84p2IHfLymckJBcHpMIboj3c3
UTYir5qaH6fAQvioc7gTiyEIW4V4sE4Ovm7VpV3L2E77eQHzSj4u4ePuxHtXxAGKJgOmZnRb91qk
Xa3aYrTXCdrTEBvz4uckcdoXFmbbUHeOCJmf7YJgpONrcBZe81X7cqe0kKB9KiLlEcCMVkr0ggvM
VldumOVp+wrcCdiKARnbJzeLDyQ1E5UZAIWm1IHTu+wEWrz9LLYpWMybgKlwy2d5+i5+j9SQxYE5
7rcLPk3HBQWDYBjYkIVc7CZ33Nv33P4ACG2T+jZ5Oc2Uu/tHeuB0+X/IT3XwENIj06Dw/8dAMvcg
3DVLuC4VwS896/eaWkPcga+j49LVHI90jzXXn5/C6TpDrdvy724tPrgWrdtUGF9DC0/65ujqVLGg
flX/x0WnXXVMvRIJhidPrX5WNvv/eO5Qy9pQCYdnNXtlAtVLZ6N41N/ZDnbveAxFJTVJVuFXNx6l
Lkx2XfGZg48PAMT+Tya6c1mRQxvWKf++XPEiRnVCwwk4M+iH4nttsHoILtCh8kkSJKT5mqyHCAnJ
7Am3Bctwrec3RMVfCz3yVlN1xJSJcb0VgISbX0ttGb0s1c4KZYzILGfzOqohhLj3/YchKqFnh2XH
Ze3EUmQyTR3uGbdk320qf51Jpx2vxBxTgjME8lN35DAfAys++QvfIq0Ipa8cYX4FU+oK6xD6hvsp
M+A51v7kn+V3pnwpEZddPXj0QBmD2eEN2v5REZgILMLSw8DB6jmsqWML4lx7uD0S6th1LBFSNTe3
ZjRg6lI09Iq690H14XKRovl3CmsbvaXIAj70AbufByr3Bruwh01gke5sSk2VlD+DbV07EVHHLXsU
UrIRm6tILtAm+5FKt+tiI+VbZBbV+9N9jm0H/s3EHgtwOLvaJgUk3hn3LAbPxQGGCcw/pTQ0i+iY
jPUL+vdRQVuBpgYiGkpbx+yifC6GhXcvEhae2qXpYwLffhYIVYqVBvsWnGdrGydToMYBXMiaX1Fz
cTXiUjsZzP01zSzeVy1KYixHyvjCDUKh1rCroU35ljR0ip+GZKxyk4qJai6eKul1sYDtfi3RvG6X
5asIcVnfqOMSFPT6x389p/Im0LRwQOhtBb8iyMrcjzCtQVY+WKjjBUXXqE0N8/gOsBTqWVRah2QI
eidqZI6Nl+NabPNO+pYK+I1z/wDv2JB9CiAvn4BxXREW6dXwNkcdEyl08IOwaKqBAfb8rTiK+tp+
mOMkJNQOjmJiqkXlbgIsc4PlBq7LiEggFjuvbOO2N9htkfn8dCg4yR5FPpQsmmgMzAqQ13x/zm2N
qKw3qJNAKyBCe/1YagDwc3fnMO6y7bp4gmWWiDa80/SrE2sL4YFmd7jO603qgw+Q4AgZQjb9fUmv
67epQ+bAJGaL7wBhlj8mpBRuBaNTEvN+gBwWKKfbrfOpR/0e20LikaDPq0t0C9TH4d68F6gSqLWK
x47qukYVbh2hy0F413/pBdDIK6lFdQ+qdHvHX6zrfDLffAQMyVOxpaBzPm5vwi1rI/UWj97dnx6v
89vaOp3vVYycoiejCIhGkQ455gctbQXb5LjWc62d2zYpEJ/e0oKA2gn6UEALK6iO1C/ivk88EvRD
oWRjwROuOE2tg1lZ9HRzleksdgyAGp1gL7wTp2FeweH5OEgI1hFngpRLfPU0ZR5jG2aZN+ENy0LY
wR/mY/plp8lUcxaD441+IuuS6yYJOG4FddNdZ7I2pid5ojy72NxvtXpRbwg3K5YxKhLcpKS8xdVD
jDyMtRzImQt17YBGGK4usEavBoQF/kbgI/jafT8d+XjNjwdSVw5fY+bbbdbEJTbXT9kMCfUW5Mqu
Icd4Hh60CIBuSwAtGSllU2Gf6MhMAIgIouXztkeOiuj7SIMIJEevXs+CqHWZnPwU0zdV1MJsxKjU
1/w63Mgsp6av8SNo/1UxE/9L6vyakTCyEvJoe1aplRiHB3AyxSfqHh5pJGHjTdBsefG5S7ZF5D5E
MN/zarwZviD2tJI0nIMhOfMEkNGTRtBKCGB1LSqw7hAXatbwhP6Dz5c1HFdIH7fhTXoxTYSL8RNU
aRkEXgm+cJQf+n7dmJZnxug+zW4rpLQXaPFdZojvieu0llGsOGTCLNF8ZlARlzChLjzGDyOs8d9b
HShqPGpcVjSGPrTJC4HRCKuoaz6mJqiHRP8ThiRi1DeZDoc3uSc1mzITLiUAdLtCRXqIYS8fIlnE
9KwJNhQx4qpuzWsYYwyQb35vqz1OQKCtaQzGN020GHx5Apr/jEQQfWRW/DYz55zOaogtd3FecPkt
Op8bojXn8HUiVw9E1ydbOfEwIB0RKdku3OYpcOXm/zbT8/S89M8FqJ4BGCKQE1zrxyHFAVT02zdX
nzOMslcr8/f17H0JKBtkCTQ+DtM1eotz9jCpLf4WP6LPlSBn0cZkGc9jgBCyrIsm9XuQ3mvRCuEw
K3f7JyU6AeGvVBqoty+EFofv/TMDOfsusUeaytAN5r88r+Dq9ZhKvMFcOX1UI0uG2tNkivqXacdF
rmVy1RO4eTfg3FHhMbsxi1cRPMEqzJYnM8GO4utyy36wSa+BIGIqMrAfqwxJE5VckKsLfLVm5aik
CzRxhZIX3g33zmA715iz70bFlquhCVKD4ybPNSzTyDpAjX5KZ6ZUU+s5/46X96UKLbL3VqxnYDfK
O3DWXMUFsQ/FcMQDTUl25Wah9Wk0K7K57y29q7l7fQC+5aAbe0zKr16h6ZD4ldxx8+Gg+vDNOjaY
XT+AiaA/ad0WTNrp9jNNfqJmj0bccdifM1RMeDFKDzwfDysRW3BeEW0DmggzT0kkU7c+ttjz+Gqk
7iGBPm0k92j6C5NEqhN6CMkcqO8e3vYhrMIvwMVoQenJCqPghxV+tetGgn2kpItTEovRRG589+cW
CjhRhHmFvSW4p7vWL8VUUDCzPnDk99ec/f1CAG76j0C3IVAls5A7MvqEjE2MnePV37T8FmtsBHT1
yEii5P+XEW3rvfYH3tL3ybXWCW1+9QESYRmUUxAejJhPXeP6LfRWZ+v09Eo6tUDRV+IgSmuP+mwV
Dj/YSS32usOJ9xaIW3IkJI43LBlxzDc1EkXq3k+M6mP03IZwWO/pDPYBwaCd5y/G1CixXKnQKVKA
uuHDyYpXie63shUIfVkZt6nZU82sHFYiEXIVBP1o9ktLhOE7wuT3PveDzSRBTrX7Rb5WEcFEpHzW
P4rjxzj/2T5iGZMIkB0TEaiC20SW89RAXcR0PLgEOsdLoKwxikufkuttvloJ2rNjH7Nf6UXNfqd0
pG+oZ0iYxEP11xm1zjrowd13t5KSqM0fG4TpHctqpj2uPXHsXTJjPf+Z16XAHXz3MuxMbK5XmZgy
g2HMQVWDdKEekYO6MLYc6+jIm+wP9PtGmatrKwUaKrnwJ7GsPM812tck2RWk1ynsGtn+SdrNEQIY
BMNDPhJm0kflN/WEHE8Dc2qByqvGhurwZa+SUKDdpGraKmKJuyvV2DHSUP3BvPrigmm6HYzcIt12
0gvt471lBLWptvic0qBdxLv9VIhD+WAnu5LVhkc2VuKB2cGMpfTXUMfu05EVm2L3PYUitIDnFL0e
y85ZUtd6KKynT/T6TlAniDmrx8Vb40yssyoATGXnRPY6Csa/7PKfzNbXjq4rNqd5xXAuikQnDHIy
u7Umf6rfP9mrTvgEHAAqobffRZCOpK8gEAhHiRO12AuNf1gm+nP339W3kYeN+eGHqhN2JeeNMHfv
zHxYrDGlRwmmGvCTGDoThnF1JcfIfneCi/6LVI8ZZ3J9VeM8SBprijDpX/HodmYppr7LeGq8jA7q
RmTg1rL/NhC/AjrtersNXzdQ8ZrDlI1Nl7m/iDn6PqYQP85S5JH4pqJAo6QbHIQ5pkhyzQKW1K0y
vMFX6VUPV3k6TNwkWPYCawBe+eFMf+1HPZOu9qiQp+yCzBt26pFQHmIzk8DohfJJWQzPTsFyzBd5
SYfNkANW7W/hSKFXI/bnSyjQWPfJ8R9OEXx4s76828vI/RVA70uHOWu1BTMNmYo0xxocwkxIRvkP
o7onfKvO6WL5y6KlVTboPZwljMx/GPiAgeAqijvW/p+QGrWZEFZJs2+2fT4mHHtKmuenNaMfqvQv
twmQZflwEQi+7ZJjYLAK9lGpzaDdsrK3ESBHcSnWD7kPcvnnKWw4fd5xkZpQVF0RC7uDqAtZdL9q
UPRxm24lhdfQPE/gJaJAyWEyIisLhsOC6bT38h4r6xuImJQB5UuoevBEB6GofNohT14q2n9B/OaL
Lqeatshorr3efEyNGk6FxtbHUgai6gcIVnSMYWwAVPf6kP6FBNdcdl4oFaozh8HfIoedDgzjrbv6
MAQCj/WIYREZjTlXtWFjo5hPF8WainUjllESeMhC0nLuYvakuaPtloTy28JhYeTEQmBlNzZXlj11
gM6AnE/XY+8bgg7b90Mm0m9wVsbjT45cRcVRHoMwYMcOrGIaazTGVRfI3OB9X0zYemypGUYhC5w1
WLvZ462gJJe2kQqbptU7/7UIyeEHPvnp451QBSsMBdh0SNssP7cpF9OT3L8OZpSKBlvNfwvsjZJ3
18RcR7bF1OHG4QAEtjWNKlyXllXoqHksutWR8YqvdA8eCrXUcuMkt4sHSX7A0CJ5B7+ysy08qU9U
szXZXgvpZ8QiT0irHn2je3vprzla+7A6O6TTxcGKR0D64L92r7sVx/bdIGUuiF9Iq5psL1HMiQnF
FzDUu/DOw4bCQyFAFCD4JE4mUYB2KszqPHnUN8AnTJ6UBLmGtnkoHzoeB4IQ0IBKm/UGWX/4Ufme
RLVO6nMhKD1/Fk+D4bj9UWOG04fTBP1Fg6BEbAroyn37v0OXAY7kubFFgKIPD7Xxul0LNwMsBdtf
oPNI8gnxaSMElTu2FqkhsJe8flP6QzwE26ArP1HRgHump24ObRQOnIZs7RXVNlS11WXqTWP2H/vT
GXm+KwRPKRm3DN4fFYl+UstAL8+JB8Kiph5tbI5hjdS1YdTLUZC5TOiMT2khB1Nu8AyAoHmdaKog
Uzg5T9ZsPvT9+50CilQo3APJB6uDp4NC/6Yyu/C5WmCSYAlcNdGQlnRF3+1UwysweUQrMr/lulig
7kKlvG5zUUCfnEAXzm4jxEealel5eBMy1xYVcIUZm4LSVMTzROq4WdUF4Coht+q3FCsdSnP9P3vZ
hvBjamtxL3pKrnrfOzCPagCfI4tn11j6iAWYu8atKNzzmqUBvpAy4WGr4HxCA7xD2h2Bo1R0Qp6Q
oHfZRiZB9RVZKofHOqmuQ+KSsEUOLsOny5Yo0niYew76Pco0f1+yLz/dTML8ITOUifDOm/aFCihf
kVgGOq0Pj5O+2xp7GxGhmWmj0Dz+12Np/lhqx9dDQchhof4Do4s2DcnOQ9UXxqWrN42aydF6T6Sl
bUMdwE/3MTfq90SpdBFCJ1CqwLwdNnhjHfGtGs5S21uABBvSghI2StE2t678RFNFsN4N4S8thXBU
k8v0jiB6RN9JrA7QxpG1VDlKs2vvGpqUKLUGo+It8QD9hCw1AO+8lsIcY2Vj43TIhYng1wxUUDcQ
5pLKlBI2/Ffy+8kikalXj15nd/V5iOC0DsUD43fObLMcF797nGozzHPnJPztpQ+qeN+zG77ChJjH
hDs0E8teo0DXlRkTLE8u9AE7hTpZA4PmirKX/TMbKSn3Kiw+cHoBQCiBL7bSLTsxQYC9Bdzb5AaA
9ealuH568duOsd9k4HzZdecvCfQPlAaLHU8W3lQHEnahdAE9HR2M2rTAKmYvGZTjjqYoRgGQI/gq
XJeKzhnrloK0h5b05FtRFbCjl4MIGD0qTMjImAym4XNTOhUMCoukQuq9FGUmP8ci8mbK5KtJgIdG
7ZFmQmECmO/S9fDa2yJPqa4LyPBfJ0xS3Xdt+citTyaJHt/ngC+YqmDlU1pFnKU5x7ZMPkY1HsWI
lfhzgG5KhdQVa95iozIBgsYR+gHHLXRZQhgDvOP1SSlk9sUcMzsI6/ZSTKqSVmECSxny6ng8nS5a
rm5mCdrj3g+Km0OU7CHVgqPdSSlm25NqgU9M5iZxjCsULTcMa28r3tKe7d77g9O0IOSQTCvXRCmt
4GrO1mVUBtxWIa/wpsb25DxlYdtyCN4/iBLhMyW5ItBgaBCji7R1JK5XB1YovTrWnPNkHIjzUcnu
c3sFztT8ZvVDDhdqZlr40gAacaFTLM2B9AIFDaX2paoThbZVqIoOT/Rmo60TjFL6b4VyYANgUhfd
WlIRot30VfJ9WritaKeJAVttRqNb4hpiorCRso77vYQMgQFkSccxYwVWLNzMQEc//RgnA0HP8RJh
BypfPfzM226B1HlWhQlMsBjFioFZE4WY5FTL3M5FuIAo7muVsEe8HaxRkOHzF4drPyxsQFoKJWVM
QcyU2MRM1jlI0vCCPntBaqrjIZY75nRpnpDLoW8MiR4wR6qw3RUm9duCOHUm5M6my8d2cnD18BWV
f77e86qSEPHG9teWKr6A97MwnpE5ricDwuuVW7somBtIYzxI0Qok9Dff9J/gs6A6vlwPpWWbyDZx
mIOx56EK6knOf0gCrGdugiD2wW4sBO+AwwTCBm4RxQobieJkZMpXfpDRM8k6WZoTVDRk6LkgKW8g
l4w2DAoHEfVsXcnZijNZMrLr4EGl4946nMq/SX26ZazByZacJmXRiKOvrZAsnLNu3AxQ11f8qZkx
Lc7IUqsf3duis+LXm26Nnt7hOV5GBNAwMwoUObkt2FB++YCXOMjnHga0oDV3mSXXxwTa4WzkTqfT
g5czKtiBpKTMjQqSHKUQ8RkOnvRNmcRUr/ZAADBWGyshBeWt47sPy0fQHETQmnV/Xi/Vs1uN353Z
A3Yn6fhG0LHJCIrZuKVzST1tQiGHoW6T3OSUbu3PYVvCH+qJyFKy6IF50LPcbIgHO6AQEA0D/9hn
OGJ4JMpQJ1lukbtjevl+uYzMjP8vmHGIx+BWoWyew1GOSKMZc7aI+qQJRvdAFa2Pc1Tz/frfkgKb
keOHO0QioPzPJbq+25vxmuHlVF2430zU+HFBvZk7NSbDPiYQNUivQeLjaIwZBCs6e6Ah3s6k1ObY
qn/KwsOKbp4jZBHdCLQ12PBFrfkqDArRxRBytfkqRwRG8j30/MMm5Ea9x/UiyIrFKUVJfKsmVBuy
tnRcRYQRyzJE9HHrkGdHnXxlIQGLK+kRaiE3SxqAb4ITKy+5KKdelRIqyH36jZXgW6t3Bz81T1dr
6IqdzQn+Wc4yy/Gn0pVnDJ1JNxovUxHDII1uHfgKyhXATMmprq7b2md/CCo+bPXq2hogaJwmo887
eLfAz8YCSufi/OmUqrg7o/4CKOYDQtGeQowFCAnhg6glpQyl0hMrrDZTdG1LQ88MRBTaI7w9pDOM
IjQuVrs2Jf11BMZF93wRg2pwPp5R6DPONAVtqdoNUI8JZhykowEvTefm2SMp1c4TfgQd6Cmt37jd
Omr7CeEji/sSMDNFexkgh0kP0NKWKTps80+79HPp5uCfS1aYqD33i4nrJH4VmwY8hwwDQJcfAYFZ
sVWM5WJkAWeFU/HHGsp3o6b/21jHbzAHFwuHGtheyBfjWw8tYNVA+iF7nGVyAiZ30uv4E76XE7tK
iYDKLh24a4vt4HmvgWwYKLc/bX5pXJKvflLGjSa7ZP/KqIgrS3w4pKTRQGsDUc7Rvg8MxeHGXPr6
2iJOSV/9l30WAvw6EnWQBYHcwQZ7H1bcxGk+QlO61Emn2HRvhPJJ5KKjnJ74P2O4DtE8p0Uhc1Qy
AXkoJ0AMJWk/fr5LjicmY/hDcaHqaAQXHofp262eBPgBy5EaLcGZdqE8VmT1zXdba218ha17LSI+
CaXWmRdZaY+Rcu1GU0DJtRmnnLomBlMDz9WXtsV1ZkudxmyWyqsED+8WZoj09OebjDlUMKo/AD3E
RcDwQv0nXOoKhXcHSkZoYAkdJgO9YeWPC2YEoRbxaNH3IZG3GQ5vZHpH8j6Wl/U8sstkCSXb8imH
4YkMC5EaAq0e3LD/NILuM5ReY+kaY00+5wiOlhWFoiCeFIu5KsTbsj8bD/fJqxM6bcRwbfmWUdzP
XhbHbXObUKjAXNH1A2ztrPfrpHkwo7UzvRDLpINDd/JJ8Ize+zIxiZwoFptuM3G3hOPt7UZFMjW7
b4oY0A2uvAovWZBEfZPIer7DLJW8N5nfMEb02748w1x9b7FEN7rCRMn61MGxefqyBXzdW6T1US80
PrZzJ0nlWvvztILlA5eqLnv+GEbjO/ldBShBiKPhSxItC61HXN1pbXz/Xf1kKW2Wy/OrHz8n2mcD
f767Hwq+Gwc5CTInPD1fOJW8pDrpG//d9hXO0H/y7+fbCokN1Aw3dovV6oPFWq8P6+Zt2uoW1U4F
j7RPw/IBQPqUcIyeRGC4lhngZnjuMK9XUFfMEP/nJmgFHW8Z+bUkCAd5NX9fimaJmQthvDYWaGZq
oFYRkwczDfLRgAl8Io11QHn6tEZUGn1DojnkwWfZK1if1T0iffwQCaWmyqTCtVijcXNg1tBk+7v3
5WkJXV+YWvdavPOWRqB6oo51R8XYyGQ7yFXCswz6nNZU7Za/r7YopsGjgKNs7wcV+U0ne+nrFdH1
zxBzJGrrOlSEAgHpDRaFIyM/J4Zfmgl9sEPro1MQg3hRjyo9mYBdWvCMpp/v740C0GYURNCj4XRn
geFG7nACixftYJfnQAicSEqq1D8sBTaYcQmqrfO6Mw9cJcn+YZ315Tv2ajw1ZVdat0wXNIA3emAd
sO6zCsLi1cYy8VR6E4xX7VEo0i3caWTaG2oEVHJ4PlCAAYgAHt+mHD0OkLdtRfruAIfRmenWzwPT
o5g944CBJl7EPvQtCymFRQ7E8S5L0kUCZDqBUQMmKHqAkgSgBs4KhESnP8HRHDc19WKGzgEs9yNp
/sHtDPBtHWcP3lP/P2pvAyW6BkU2E9i8wBUw8guYCJfTTP5siSv+qSqr8nq6CD9HEHGpHHIJw9+a
hE9OBFgzrtnPj+4bCzNRTLBcIGHLbg2JhtUxREbDkmcFlDgNlt62CHr39EqQ/swfk4DVs2XlBers
h+FnVoQkObj9pO/0QnRbKudy2AtXNDPq8rM6VV3ht25HZgGVxwxqlHPH634YutKHGev3KBgGnwwA
mfVi+2il94OruoAU3jjdKBWL9bYtNC5iUPtxjKltbMaysDPCEy2SUC5BeDpXnOBy+lYinCcYqVJ6
bpcZpBHtfwFVTOV/CB8YNeK7lfpZHwYtTdUFuoOIfaEs1Ip3V2v0MNGOmwY3ukibEx4/Zs1pWWVJ
EYKoUSEQkHwiFFWWPOwu608oHiAhjCIE+cQ4Ku3rSTWQH6xQWbo1eSH3fjjUI+6iiwwZdKMFACVx
YUQpNnIiiXB+ZjrupecJWpLuz/rA/MeTaJC49SRzPumr7wbOb0ufk4R6qTMjvMJMu1Ujpi9WgJfK
JzDvhI1Z4dxmCxXnZtvN8326ax1Y5joDzv3N/50dqsvfvRwM5FPVoxFuq8VGJzf/uK9FQvF6Qb02
HzsSXwoJANBrW3nQXXu2BBMt3m4MWiq/U/vwR/xYe8wJgCKkFlc5Ui3r4+okwZ/VLLgjO3KpL2AY
LfnlfKl5wyMEG7Bq52BZUgCsrP521JO0/T7WsDyiio5cBYXMcalZxC0o4D0kgdi4msTMHg2nbbU2
VCqWvJqKYCTM9n72u08QLI/UI+mrw3jt0v7sORBryr29im7TNKk7GsqWE1wsVD1x0Qd5OtkMbJ08
VQjdosW9pnsLYRNQo67iW4qEIjf29advryfUd9lHLqXzsVWfpkxfKjmvJEsyMMc/1RaNtha+e2Gt
3EgJIW52tS2NqqhNUgHOSxtTYL9DAz1mG3StMuYY613a1tSqv0J8RL4hsFc4rkfZkMTm+tfwnTXR
qrsD1crwhAi/mf/L6Gw5hYLJ/HZYGdnM8etGLS4ARkQGpWOs+hIuk8TCEZm5BQE5TH6IXbi+kZsW
O3ipr2qNC9m+qassoHUTwvDcZavykkwfdjqNHOb48pv7a46c29XGKFtln8Ik0RXmxLMGz7b7v+4a
0J/2jMha3oRySSlHzreHIOp8o2XF5WUmNtufSF0gZ4f7JtqQCwmjyjCn6UHFpGUeXmOfxdWJY1sj
FSdhAvsnCZQ8pdYXlYFxYKrlb3JvBnJLAILDNihbHlvsyNdPMgVD7SRzQ+yv8zeXaJgOYVlavPk2
4uqIJwnMZ00D01tCzACUnvXmy1sMHx9tS9GiXa2RuHxFSr11EV2/eVF02x9OUiOxq+KvelJpjrOJ
7tQ0VZpe64RVespYjFysuz+c54IrPPnAj5psmPljCuh/38ITlsBwAq325fXOJVCEfHPOZF0vj+wp
Q7hgVHh7/mXomtgFU/b7rQVn3QX8FO1Uxzwup/ieTGegYyr61EO+UgbazzUx/1UR5PaHiOw0Rg8s
liVjObisRelSbHJqxnNWOn/9cjzkd0rwEWmrkUx8I/T+hj4xXHqbASHHyzPk0tr9VXO/1p4rQKIT
gn78ELoIDA4SgZGSzLlORs2oQixXj4Gap4MZWQckL9gUr+DOSSq+r0201y8v2rJzv3//HLGYlU89
LiXR4U7UNQXvCiEzdewsb234iZeZ5OMv3pZ4IDlEd+PGf1ueE507n1f82Mnt1ORaZwb84dyB3yRy
1Qdr0FRe+4hg5R9iBgglZUrJPjidpZX0tTL1h44tE80jmJD2mDhgk+TMRWEG02ArNOid1VL6wBXd
W9HV17n78hxK0ChbQh9LIw6NXb2j4jfHoUBfgs5Wm8nIWiP9cATzurJI65SSHwVrMkxIEoyOzuXa
/FKMc1h/VPh73uazyPurnOZdIeniSfwgc3bZdzLL82CC6Wp/nvBAeWZJhMAx6mMiZHzf9xxzdkAW
u+GzY78CfywxkpxxSgw5fUD2Z1El9GiuYSpqGEe2horp5kb5xthS3ykfFFJgHsUg+x31GVsGFM5P
PR0ma0t8Eaw630IHmGG/Rj5wwEu3EfInEiyCFR+jI2qsM4iby1pbl0sx60j1Wrg1dW3QpIBUR5r2
M2uTvGWeEZ5pY/ZXdBevH1Mwt9t03zms80UgDMzT3WssaB09o+A5w2/CJeLzUePN8R2/Ay1qjssU
9AXzvzZiEya6aENfd754/DU734NHi7TLfpVaM++/xJnEmuKRVm2717aPZk2/FQT2L1cpGHeOAcV8
OaNdcw1SAssm3QceD4NhBqZsgNfRSwzM/mthN7MIssV7Wdp6ojQwKjTM5zPMPYcdRhecdZo3WfFc
eKSFe0Xq3DnD2LCnY3293rYqitFOJR7lKJQXKqh2nh6W1RpakxwoXfp+rEhoEIEwVHnhV4Fqj3rs
aHFWPfErdlxu6sxSUO98xh4gS+0ISC0oAG8MRQfTnI+6nnQQ7A7SWBguprb892/9ZYxkD9J9UECA
kslVob/YE+/i4Okqi5Yr2oWNS7vVUl2xnBRJyg/kjsxMVQciGPkoJkHnRWo77nG1wTyp0FfehF1Y
+1J82tUWedvK3v7BN5R2l8IZyltHd0XaSawlr8fgFv3hYyrRaQAU3R5XI7hP4LFZVquQaFRLFKPD
U4M0ybpFl76v9KaWnlmX09eWmRx2UMcVR8q1FydsQD6iPAFaRDxN3I0Idq/1NTm/X7eMlOGPCjhf
ZFkE67N4CIs56Htne3kY+v0aOHr1G+PHoF6JEJPDaMIvNTiq1q3Og4isC1AAnm9/VT/dpDsSLMIm
BLDQmGalP9U8/YaeLqV7AUgb8YnjfB7owi8y4OciykxGKiOT6o8n23co4INgMmzAv8t+Fs1n+IQw
kIsYof/foV7wF5Z3lSvyegS2xjVw43a6BnF9fmoZ7CChHL7nWeBe8dI+PZSr3pMXk+ivntAMLPev
RxlqM8mi/iES4oVObPvf/DkztUZYpAGEpQFpnbtS7Yg8y6BqA2BrjH47BPK3kx2aCwU08MLnjv7K
sR16bVHBND6FxzmTKNuB/dsCcfHO5FTItqdMwzSq2DBwAiYFRIH7YYKakfZDgEQ6XlNvX9f5macS
Rff4SLQY56ieN9e+txPJICwAhqixU4AcwL9EUi7lndrxmukEvxae77AkXnVfbt6jkyIxSpqnuZsO
aSft22KKj4wGQ1u3zjyycTgvXwhkXLFouQkrDXkjKwlGQM/3zbv7K8RxRtuC5iiKmn4Vtahrn8VY
iWlzK9aBgkTSit5ojxsSnOhl6ZemTAiNFEYE/+adf5KDGJ0lwFtPbjEc6Vqt0Q5XZlJhElmSREIN
1NZ+oJADyqmVU54L7I68PwZw1/Wg777Vi/sbReca4T8bOZ1kWGuY3UDMGuvJXpoViTS42wgJqEaC
G707ovYL1mkuW2ZXN6YRBteE+k1tQvyHIEdDWCTW1ct12rVbloSHWroLxZCYBgQz3sv9YDCqWgow
UyOzc+x/HjkMHzH3Ow37tc1KIL2NzNy2KqxJxXzH3sHgzZznNh5wG1vlz5vUANzGlPAX7Ls0yoFo
icAYlZO5hZ5onFfN4HLh+7cfbPxU4U+KzkRPLXOZ8J7cEmz+bOdmmbZfrLckoW+qZDQrpmQNZXMs
EZ4mF+8JXYFPOg1oon8LTeWkNEkwkunRGIKm9j4me4HSWzU2RDNnawxuPsC/zFOcblrY4tPNt+eM
xpNdpQJW5J+oLkXeAwFiQs8maoLH/zlLlO9nXfklwRnnnI/qMeH7hymkP/RbcW3GERfJhkVg59tI
SrTTHMBQRdiuD4mKfXQdS3MkoD3fCWjkYDlkAimdggqnRbWcLoBfkFym2VhV63xHhtTYakJbBqiX
tcwxR+QhoGSqW7xsJmwuxcesEQE2Fh0iO166iZYJ5QKeM8B6czlejPGy5YV2Sr4ELXVfP8QH0/xi
5gROiej9m5q8zrQ96s5HYs4HU/fZiUO227YIGncvAxqdxv5ivxKqa2cmUdqAdEOaax6+nSdxecw3
c571+cQc4onWzfeGyelnYsJYc+EgOYf1VTrtfu8o08bcFe5i4sjEvCG1Su6TYYieqnYXSn5I+qhx
/3FeW8XVojB6xiawUSCnb/+r6y0CiL7vgOtm1A55hZ+4y/IPNlgACBuKyALTxlr/2FxPLMhLKizV
qU6icHEd/T3xlHY5UDtOEUduQ7YoJtp+NFyTYdSi2Py3TFHx01NMNXZIENlTedhLe1PLAwTMQFzV
LGk+0ZEJR2s5oHkJR7wOHgdwEL+2uIiI4r214iaFSuJ2r7+0BGjz40S3G7xfdSZ4JlDf4h2JFFsi
6k8HhNFBVRGxCdjtbX0lstE/Aoop+vemyrVV111eVxjK9XEV47DzkDQNsZYcaIy25IGS7AQNNSoP
ec/8KksLSM/bOPf/+OCXwGuCnusko8VfHdRxeZviDJ/04aydp10Ul2hTNh4kLJ41yRFF/QuHah+k
cW3wkHF2Ot9UObjMBN330G+k6rSgB68kJa8GKDUUZ9iE7gDVdQnm79AvYz1OdgAh9Qr0zoxttvh8
j1X3qKvLvOr1lq4IJnSCG/SAOpLx4T0pjJyMRBCKaXIRdMZcjrtAJzigKpmgplYLuvrhk1MxxHS4
hgoOFRElB8IfRtkuW2Qv8Wox01H7wOlx7OprfwFN0GzOpMgRDaQeg9SVALfYf+3j7+rua86gIUt5
6Qz4oaMBzIS72HlD4N0VgAyHzRjOs7ffG4LCf6fT2LW19xuehEfXWm+EqgdC2MR3qkef9wqmir4D
iNlIM0sXpceiEMfcNk9Z0WjSniqiYzo9rIDg/VRRn01v4HBmwVzpLl8zI3yscd+Tr0NkVh+YFrT4
YivZEnJYz3jKu3ztMwf/ekomEwG/7GGTIUQEaaNoi/MMJbgCjFTOcUu1JhOl76hLfHkxWUD0fvSj
+qZSJNp/G6yCsNatZQn/Om1Eo12B+lrKSPjSICHcO22eEawM0Pb22eYtbxuAU+HKPYHQrI+P/+qB
WlMOTg+g33jjGQ5Tv0f21LZMfbekGXOFm2ViQ+VALd2YM4mxpOVpRzOmvGxzFJwkNv4bbMhSLJaI
6fdfiyRIJxbLmlpgw08BhSodIJRBzR7fupSX4TOQ//yssqpLGoNw8mEjXXbaNRy5sq3w3y3CE3jE
mXV30ngZO7Ti/Z+9IhbP6we3RwYqVSR1G1gb/I9W0d3W7GYDZ7i/WucRct0T8K4kr7J5YSKSRG33
aquvMbsj/Gb+m6KN8EdxtesJqIPRVzF8yUg69qeycLpzzqee7S+NgG+ltnx7J2d3aqPiKuaVXVdZ
uazH/AmFEpGknKoFLH3aXPYvI6F6+73XZWbCAUT9wzfXyGA0LEw3d6LigdpXXeVTLArXMDAQAKQw
dfapZpV+Zv02NthOHBfv2uIOrCXoh1He7vSi1tRHNsk9PVRS62nyybPPum5svRgOuSicdODw8cXg
HIydz+nnMllvHvOb+mbZYPXBoIz72eGPqbHVNCzCMQxdp5LaYgchiLZg892p45wape6NT5LKtAgL
2dJqF7p2+dovBQgjTDmSciXjSQ1zr3nLsYIVIL8HYfAF6sFNmr429NJHCeF4dQ3Vm70QPUlN4duC
zxjMCwPSZ8oltcxVruF76ZkecSJEsLzxBj2mGxQviPMkhMLIsqn81LDHGkTWiRgZN/WJ2FPsOmO0
2Hyt7v9thJAn3FTIqbF7lNm06BeFth5IcDaFq6OxXPR0ZPxcBE/z4QQeAkHtLHeYoBYfyOSOEYi+
6eQg56YPZCb1Qlgr+SLXS8ANQA48D2yBWKERvmG7nIDCOBgpdrD5S08vuPrmXcAxHknLUERuM3K1
GeD1noB3g+CZfABkrOmLzUfaUU5OHtF6Liz5jMeScAlEBRzzlr8SmdjwAnyrP0FG/Vj9g+B9ogCO
Z4oZBavGq7dx2sweKtN1DEc1heHX9kdG6qSOZ3ow/16AKFX7BAYk6K/x24RiNr8qPKT/UBS5Tk91
joHuhI97BpKwTyYDYZBIOEF5aCuoI5an63iunyoPrbyEHpDWfElcPe5Lfj1IYhQhWZUgOiP+6TFU
dJO5fxoXVIUJ0gf7fIDyOgwyHv4+x2v/xQC6D22HIpgmkDYlfBXnTyZ35ZnHJ7veHwHU2SSGPKpU
JHn06RU7osVQh9QY4dBWioCorSBhAEr9pPvzb0aegFG9wzArXTQ6kobkAHX9BYP5nDw706IOfrZA
q3zR0bSLlNJoES4BdfQf1mop2eO7UmlRFe6MWysuNGujoYmAhgWZJayNQJhaA8mHSgwkIOZTbOoV
4/gXPlYN+qCie1TqveHGmN+8wO1Offe+N2+ujuJk4M+TdEyuPO+6fSvSttwI9QYRmQtOd1IaP+iZ
Np9+uHJKZh35qTBsiBj5Brs9Ca5I3WHp8obdm0qPLWXENI4x4IuUY9/KC1hsN5CKzGiGPAd8lriB
MmpkhQL8bOjxkuI0s4Rrp83QRdmQjXxRh5P9ak99Ysh6WijH5f4mCsQQL4oa/IWTpEYIR+RV8qZS
PrzuBkGASUomEokTQitWlwpRoHGeu1HfvU5KTOoE+fzfuzNfBCT0Fdm4oOBQwWGqHsP6pIAgUhG8
8wab6P3+eB9nkn7x2k0oLyhEpekixfPFjpeX2ApyebY+p6lL1AvAFBxKOzGQkI+F9PLzSG81Esia
Da/CDYY0f/YL+MZWu0w4vQqoA0ysxXgP6YiSdy6KgF9WRteveTz6izWLLjlij9wtj6JnNQ3+Pedl
96JzG+TafcEZqKiq4FbZOaUlrNfMqDQjg3u0tSk9mC6xIw1hqQmnMe6zHRIs73anW7g8wRmwuj2G
PCSvWM2CVld3V20CYZjvS0Z+v0dTWQ78xpwlFtmspT1YP8uwba6bDOaITjYg09gohpnLv5rV9O4R
L3iEWog8yZd89vewki+t8ocQeZSpE/ZliiIiB9Nctozb//oMulWZWZNT2rwqPa8F5w+1fk/TNT71
yH0l9gSTLH24L4pLsU0pXvGAkg7L83EtMknqD5NNpEoVN7nLEoYJyh0dV+aXL7NU1z8VWIaY+R+4
UmBttTcadkBXEVSwYDXVYV8u+camd+UvdkyYBFbRpwVBvdMnQLuITDniaRIExwKh5LdDck7MvNoN
mZpcpGjuwjCSbdWNbuuXHY5QQ28JnAjy5yVhsAhXPmYHz78SyqdwvWtrr6LV9Ewzp/UDvwvC2tYF
/WWV3dCnYKaCCqeFpBMPBDGcb35b8B+CAb1rN3XTfcOOS471KhX3zdfUlOcqZlatD/G+/b1Miz9f
tBn3JXf+okBcdQBedpORasSCIr3Puk1YC+Cb8N9iXSPTsbl/vGd6ESFIRKgBuCMW9cRwgEjig+Q+
sglPmBWYqf04+as94jiOhtXjmBnXV4lC/wAw3tc+ANe7tOZsTUb9CDM/L4JOZjDGkXv/R8gmNz9/
zDwwLTSj0q4XHMJLyNaFHwlsSyGUB99lTb04RfWBMkivEDY8OgzCTBPgrOdv/PDaeQZFO6Vp0qyG
J0jjUcAz04SVp8ofDmMTOV4G81M0CSqCIdkEpc/z55hHz2kgqgpFywXXvcz0pwfM1t41MlSHTvdv
O20H71dhgLjKEu5NRcCtRIbzdlBDoh1KOdS/T+lEKztV/WkHHgnxH5MxAe/YEXwPHlZTRtB2zJ8E
eQU2m3LRRnqwMvcRJzqrHI5wpNJFcwQR/ZhmUjSHcIF4UXu7usEF9oSxFdHOW6uiOHGcohb5iL3J
91jXnlHq1CGml+vfEyhCEkm+bH0i2Ti6Lht/6q4eLDCuFFdTPvlM6KYFqB5lULawe6zmZc5huA0W
9dxlNqGXig1aqWwMSJ3WCA5IbUa4g9BCi648gBOkZ7l99y3wvCAF5XkqxBSjV5Cnq20EGFTkqUku
epS2dq5+R2U6/TiQDPaV6qS3MKzMTPmdYhGHpfuGquDCsmMEZkgA9KRACkeZipRH8cMRjQhhC3rD
9avCM9johH+9msgQ/XAPYSF1eIaRXzugDSCtu4tJUbVClUTEByIIiMwC6qT0Ka/FR7D2LtRRwNf1
FDAkJ8B4NlunBh7afgs1L5VPc6wqnODPwC5gyhYxSw8MR0Lax2bJ58dIf+BAovwWk9N3iLyVjzkf
Jp4rmf765NIlrLdomOvpfkkL8D/u0fUoCZ8LPxJnaSqVxgu57+CblNENQC/sMlqr7WafGl9HVcmK
MfpgnMwpfgiBbiUufkBu04ABjuC1dzyJglhnv1LOAJobK1G9Z2v0ylY98dQIz0rk+jZcZCB1FAqT
OE/HL6EVnc3TRaLBbXqEdahjjmrBGdM+0rv7njRHDpTU91EJXcO983Z2VImm1G/ilciBl/9tC3UC
eTokyz792JuJdW0CpKvwJm0bcKujecadkam/V0gQ4LKBvl0OBC/tvGeu0ntF3RUBpxSZiDczRiM2
8LePO/3Gd+94plLZULNGWWKxDzCOqwTFMIT1RXua4l9B8951bvbxK2q3CTArJOiR2RRucLa1Gerc
5eAHKC1Q1tAQtwlOAQpa/aArJNXkTjWj3dh8JnY1JEYSbRwbIx2wlVJTciEKhNQzsDNU4BlFEJyz
RqPRjlnemwHZGN1nSDGOdsk/jsuZ+/vRj/zEypW/AA3eVjY1NUK+qC1a22ImTUvRS7C2YGima3rc
FGjscv1hdV94fCcB4O8dUdxTj6CRuoqm0o6XkdQQfT2hG3TIe+qrPnmUvbRCZf/WRd4wVq/HOSLt
KieXs+Pr9J/yw5QJSulyuZkY89O7StqZKxw2yUECb6jIc82ji85sKBRTlqs4YaF6BYcowwmhz868
D/08aSZYySKS8CsDORSX+uuHScbS4zDwVKS4P2XQDgllHmiuDisJh45QL+tYwBZ/jaGt1X19KNmM
egvDe1yJRiAS8QRbg7CZmq9GPp6sY8fg3FpcU0K+T/GE7dth7XUEYnxNIlydqG2ZP5EiIMKK0YJw
Lvv5IHpoPLmNc99cs+u2dA8eig0CaskBl3cg/Vh/nJ1+GvV1kBsKHl5dJROLZ4GC8UHNIX9dUEcY
SzIlSp8N+WO1AuWh5bLeQCAuFeLvo/L2+GZLPgt5bT9EM8Zvg48MYODyVNGvDmuHyX9EUKhdL3l5
0/rgvzIQGeg9ClbrbHy8ETsOk5q9XrKOPBq59gMNpKjaT449zK0qCAVeC2M5PmtKMKCzR3HNIL3+
hKhAqD5ioQONk1KQbt0xbFkFLmEmPMvjqz22T/paNa/zSbR/FTpUu2UXGpFX0XUu8pD2A6lCRHcN
CciFqPVdUgneXxLwxzCewXoAs2nRyRmOmnPpgNIhDSST4hxUSM/HtCdabQTahfFdw0a+NkFBRzmk
udFGYolc0vcBo2B+XYb0imMFughUILjvUsNaC3X08MFKsD3XpEB3M4iu5F9y52f8wkoJIOINxI7b
nDLP4zTAC97me+eM5GD/qmaBg6UYEqYfi1GCNyxNUlkmVtBYIuE0y25Xyt8JOGBSMOCMdR93oiEz
TvQOb3sLoefoExHT/8TRH+xpwjAP9pkdO2Dh2kfhrI/CdsXG1zcbf/54TRKsOopHCiQDPdiFQ1h1
HkQjHtCTjbStvWOL0odS2MjJGFX9uahQYlKGmOScauStiMw/FbmLSRmlXUnFXZW1NSPSy2mq/jE+
vAlvxpa9P8TPPsrZg+7DiNT4iV6j4Z4TlaWkm4vSv+b0hG7N1492BjuYeWV+Mjjh5WPyxGZqrgd/
6QL4ErjEVPznbfOP+IBu37hWrrEurqRX8UZrIHN2UCYh7AOE12+5oFAdo9Y9v/Muhe08US/dMP1g
v61SvuYRAyKmNZUBhqW+s2jjf4A0Skj0dMO6X2WZWAOYlyn5VYtTthnjlJq7upJkCshrtLFw6Bud
VS6OaKGMYJvvswtLdejPilncJSSK7ARtMyr5Pao8A8LZgr3PLg6nabtAGvDU0tszD//i2oe8NX2s
xCo13l+wQBS5IOudzlv3kXRhEZfh0HSW0pzsSljMgP5aY6uQmx1KPG2fsyWbOMITplEjsNtD0DQy
ts5jmW6ZQsrmDU/OjeC/lZ+nBGZZ2ZNfraxlpgngkZE/Ma8YQeabrr0wZV5A3LDgXVmbtiY93fjN
Ggh//J0BpFadbyhXZs6HFHu/dKUfAcMt81zLIPU61kKWs7k4Mzz94u8qIAdHN8MvACGnk4a3fwDT
7IzC2HZpGvISjKjSHAh/xFt/5TXmXMyyMFOmzD9m2+fh4y+VPtwdqCcwnDULTDvXShxU4FTRJ9BU
A4NmIvNrlRDiOziAT7puWW5UPMhBaaXZp1yA4KInKn3CVJ29WuZ2CW9lK6muZyouhNrueF9jyANk
q2TNSkX2F1dAPZGsBM6uE/9LPYxnYOfB1HhY1M7TAmCdwY+e1/q1IV5osz8Ay/vmGhR9QVaw07ZV
hQnlvPpUlm7Y7/Xn4vgZbwpw5IISROG1DjGsGaZKywETalh+oOzApBXVESPv3Oh5eyawa8VNeT32
eAnBjkRgg1efjGU/zjGu2K0pUoqf9sjeF9T6jDh8IAS3VtFG760lzBmhQxxNScPUBc9CsBdFNz7R
Eqoq4SWEe9isGUAJKjPvu65oKcyxkQcM7tSBr4chNcIrfhhq0j7lWKavAZkkvbmaOR06U0TouFeA
9mGspk/ituvEqYG9G4cjMCK0PYaCL+SRF112JwYrw7gShktr/7RwNS6sMudD2uZpzV7RaQkJH24w
1th2Qb9GfTLrVbo7xoHsaoG9kK+TZ38CHhhCAXwkOF0re30i0MhH4J2pbNT8YHwPi5Us1G4kSLaw
eLI4BqxJs9/nzGDUYm+NMzWumZ7aV4TXITLfGYaWxtXR5Fwdo+MIXVfrq2AGZiD6JZ6LThg8W/P+
9PT/8AcKS1f5sFFe17eHotCHNdPAD7oLmaEEe6TtH1OCZilL0XYKMeREBkbc48mRVi+NFSrP99zE
SUjm8cYliOOS1pc92EASa/d0A7x/HSE/fItCPvZf0M95IiI1GAGpG2z9kXaQyfeJlj1DGihwcyzE
ckf4+X+1WFSK5/eJx+uqpaCtq/hkihvHks6rF6SsnYDbbM0rqFMxbnhekWBXSofGtGAffzPSGtJB
f+F9HqTqGpC+Sn6gd0vSz6fbj3U97AjvJtR6h4ADKqU7+7zQjkemUKJj2RFsfguscSZDRN52LDyk
v51Uq2sZWaM1PRy7d5QEQNv3qjigqyly53OuBWybgqMu7EIkcM8iup4XUuu2mnysks8rNwb7Egej
52uhqlGaVLT7Y7EwIj4qwGEkdSzPuY9VfRF4+/fJbZWgeIO1joNNPWXvx837b2ScSoxGp7T66+9o
2NcNOgt6uOq5P3H33HsfKgrbyi6k6jGhUYXePCvCV7wdcyDGvcsAhO+7ZbTqeaIcLdVy3XDzMNea
Z+cNdWZpu6uii1VisPZPvyLM5jjjt1Hsv2Pk38P/ojyGExk2Mtu7U2x6U7eB2k/eHU6qqBPhG9m6
h93i2M2/2ej3yYzVK9pJlnGUQ7ownMBFcv0/F158RuEucp3mOtV76fU+i4KaESiusuitOPrsfEyC
eJlWghUj14ivKtdiRGAmGy5U54HxTTwi2g4QVDV0zgMe3yAtjpLH70VbbZX2SwVCIT8CmlQzsYya
jIBxhV7t3/0AItpEArY2QhxpQuIpg1B7UzORwSzjx8IQspVaqwuacaCGwo3VHGERQTMYXiz/eMQx
PkfictBV/qNLw6Xl7sJa2sCRKmkfkb4MELX8RLUPdaKqDr3yl3wdbK9qALay0XuSxrCRirLzDbYv
xO/KbsuF4j8+qJbfNTh+nvY34Y8rCiwq85o/pxMQ8cUhjG5JqLEKEXOcaolTYKnYqYrSPpcFY91K
VUyzShhXPllcUt4VP7ojXqAAF33BOEHJxhzHLHdy2qR1XE49DJ4nkBcrELYVxHe2apMmRHUVkJSW
VIN/0PriVD7jHycsT77f5MLCShKAeSkIM6mq8ywowExx0o/55+x8aE0GSK+3TrAGldWujsDIORA2
8OOm2raTCcqoJvDps9pLghkkIAruz2b0mBoZyvYSd36LcNdNbQlIChh4RZSZfipSbS8PIxBHd1k4
WG+jCBa8f7Vd5Tvj/WUHPph7yZnZu0+ilBynnBHH93qdC4f0McBZQCz14A9o34XD/ls4m1fe3Vu5
e7/MkOU5yHeZv1wVL4dJJRwu/JPPGmrNdCA8XEqSaDgSZDjRuhhTl8TR9pYpjkrkIIkg7AeLf5eR
OJk3rj2eA2H7QW6Rpor7u2WftA8OZ4Sn0cIDErYpilOKTNoyt/Py7omP3+J3V5OiKgKkyECXj9k7
SAtI+0qVV7JNq1b0XjP0vM6l/xGmAhTtd/5JFlWoj2jMFgyP53KAiKAoQpzbkRM4x1SGNQkPe9i/
VyRY0S/6QAi99UBiif6i+kV0fou5xqpeD1bdxJ1AGrSjcjlU/5zCPw80MzaNFmfABFmnya7ECTM3
44tgkOvAhkUdScwiLVBXiOYcQTKtGrtLzGntqYXg4RYC+ef/Rbije9SJb1FE+e3arL5soNXn0jAR
NYWvJ0GIYZefZQL1ureVVu/Yq4MKpWh86Cmg/n03GnDYDarfM/jwoPbm+qmtXr7frwyo+hKAZ2xH
c64cZSJawzhK61iuBJi58YKATrziuhgdKWw+294OCE+9v4mHFHlHAY9SpJeR6bAvFzKERoBkKNxg
gJNpL5WMytDalneTmfMRffP8htwMrwMqZEHg2ZD/jtNLFaHDUxxvWkPBFyOkXBwiOBJ7cE0FlZ4k
PnYfi9EY5B9e+W9bzrOOj58XITuDE4kBZ15Y7iXkItppzMU0AS6M1NuYNHZiRaRSIwLYXKNc+4UC
URpTl0gj1hEcYU+IORGdeIJy57CK5/hUDvkhXR3qb4ugH4cn/JBf/pveuMchAcR07HIpUK+V5xtl
98t6xQx8LBu0MnYdjFJCqOx3P/WR5LPpEVr/IPgpNbw5T6/CPKbQvUvsAAANEKHtb0LTmyOAabfU
vyksjn9yPowQWF8XBtHlFiIveXrEu7dk/ShzLVtZpf3S82VFi0C8gXwn283lNLemfflJycRi4xzJ
HzgNiG6lbB8wQl2LbIgmOmPTmeE8BAhFntVkgx/joTicKcMblBb6phJoLWI8psmq2IqJ7wS/kH2z
qbFtxqqCs/0HO1+k0W8GI+Nfua3eMnVR89c2v8CE9rAY9HLNJW2+67fyiTuwp0jpHC+zc73RsijC
E2YKmEQAu7HsZblyavafRg7+ixI00g3UQ32Y89rjNmdBmW8/jOllMW5/eBQIR84GdgsAGH35WON+
CFuecjCtF18pp24DgE3zIGTQjvLH1VZ38MdAEJj7OWBdW7C1toSxQJwCBXJwbdccCRApEwlewYPE
JAp+kiSr43UFVuuL1WQ7oFYuZP7PRZL5y7yx0NvY7uKrXmsPYP3gqNYJT2DsDHtIGcQlXdxbMVqn
iTng3L+8Wv1Jbi2PDZ9856lEvpWAz8z+TtB8o/qm7Eb/Cl6lGfJsmfaxRz2Vs/igzA2Q3IADqLQG
YqGBIu6p4N69Tg9mPFmA7mmB1FAGNphM/lzZt+JTCA37o+UajQikyVVSzNcbzbvNsPlSIITgjOBV
9UJUsICknzDZeIzDrAR3Oaxp2hAj568AJT77t+kS8cN+k2T0l/ysWmGtWxYy4mHe87Wt3EqB/dms
R3zwg5yNB3cOyyAH0yOljCsvPLoJU+d18oPmB61vktF73Gn3+kcm7e4POD4reHQ7L98tHtOV7459
Qkdk6NJ9s42asQKn1mChXdj9Y7Y4l9NQNCRsJpP4oC9fiOvZ8ZUNkrFGiKeOKAdh9yFxRhRfSLGr
5bpXLAeeR5xgokIouY8vu0YLRDMITjL78xH1kopPWJ870pZIpnGJ9BK1H/jX7SNgABrKPEVWS0zI
Bwku/tjtWwkrUzyk+DIlv/XX8cxi+hDHmCYcQLkdp/Lj/pwRJpCZl/cgjRFd+Y2qzoE++CQcqz/X
PtCcu0DUB1kcgqHie2COs/Zy8FU60Z2zK2Dhdlmk/FKHKL212VyxePhxEq+F/04Bosa8xhxIqqjc
3nBlu2cPcuNHDiIEWlWb7dAW1VhpNd3G2SmRdnU7wQZCfDv5bPk52gkTnZaFqqRRKcc3CZxCP8IF
KujyCx4zaVby4v/H/dTiPh01ciujPqf/KLRUoQOJ1KH3EYtmUvGnc6tVD6Rai4jFcdgTgpAOV6Ee
z5mlz+EIMdFg1lN5e+qfU5BnHUBq27ILUX5RCwY8aBy1xlOEIEPwDH1vujIDNUvEQHtgXEawD1hX
KZ3zR+7K+0KdrE2GDxY0PWoUxbpd7ZannAQiSx/XVNUJQUQ5S9PlVwYTbST1Rnd5whwQOqb4O33h
IJy6AB6KnF5a2G2/kk7L/bSQRNwJdyakif5uHdTVnU9H5Z3Fx0ea+e4Fbkkcn9rC3sLiqyemplzX
1eGzPH+77RGa6SlxK46rfPrqUpbquy4SQaY90nkMAvw9NNQ11Pwk7FQGPkkm10CloxRQXC8tJvAa
HVhGl4AryKqP93+v7DzdiPo3V3mjrhNmXlKIy6nuS0+/EcYCFmc54bP0g47gjh9k30awkOACSsg1
5/Zz6EBojnJyg5QH03eC1LlR5D9cZPdEdsZ4qXIE0GXhnMDqrPxUafPDX0gsgWRzHYVWeLrXvSsI
0iJkjDv3CBsVYjnyj1ldW9GSKM11SVZxw2NnZxW0gh/tJGC9soK5Ep6T1jN+CVaSC9x49PA1EElA
4zMFdySacpez8gzT1tBjyFW5uRTGHkJSrceNXgMPi3Chp3TqgX3uv5ZslI4qUXg4UkgOycOnqcnp
X0U705BKMF7cHUdg86UttUzPy1F/Z3XpnFVxVDVkTE6J72OJLMxuZYGMiSdKpgNGnwkH2kF30gq0
yUs80k1osWdiATJiXz6nsncKYLmy+n3VqRftOmhLYBvVWcN/z/Yu0sgU9j0CbHpvXpaTR5bVOx9T
3ehB9vad1ut6bf9OX5QWxT3bphQwd3K7LTWyYfy932QqWz8+eC9k22uLnnQZCF337vCvHUUDlNxy
5uNpZo25Fnb4eQ6hY4Crg+qrml18Eyou4HmBw88CoIMf8Bc2G5ATIq0XJfD/58vA1IzFEurfO1o9
atNf4dRiUOs+6xVBGLUXTVqEgkWt+mkH8nClf4zoAB9bih0SnLs8Y3k7AKMfNdyDGO0G5M7IUagw
FO7ovBFcTRDD6j8Ku9ZtWt51fzwq9wgJqcQjJegvHu6K+LVhsmBxqbaQpxRjBKRhTxkBQtaitbfB
tVqje/hAbiHC6yhLn9frDKRT8hstVL3dhW0yOkfvxokFVQAlygT93hp5lu8FQf2Xt8W1cME1oyEW
dQ2DQykuSoERY5M0BOxaa8lxwdIqi4osz1nJIclLXouiLRcD7Rz4E3d/x2OwEmZpbXIC9zvqH5W+
IEjsk+UQInxMnahcTz+wg7McV302YEBdk7hK0hBLMAsWwBzXqPrb76yDu5QcUB66xhc075j4l+lU
R9Pjli78v1joOqsjeg7nfwFeHaebUoBvYDeqD2onsDXXBbYAbXkMabY1ouhwn08tfQPgtbVASeE5
yunDkKyTt8K8SlEkwdn307i+7KqKgpYOTjU4vfSG4hLISNt3yYXwIEVUQ8dIfuuCwvr/W0sts4Pe
gnNQrqnIMqw9NrGlW9458TEJvwnKhZPPO+kxAoAQ81Rpb/T8S+K1cVGred0NciQx4lY1J+U/wTNi
8Co8Sq0kuzVCR66axHaJjoXUCSOD6F1HbLDX8bfPki+c2B5W/BQFJOpmCsb/lZYMsF/u3z9cE4YD
SXIrsyhkonibcN4vuhlkc3SBVf5a2fc47bN2QNnCb/qSNCSd3mEu8Wd3yPEBrLp07WWM6/c2NveP
CEN85H/JUFrVlT/No2x6z0AWPv59oX2HlCVsGebfiDBEaAiQrMTUlgiBxv0qWppxJsmakNSvWADK
Gt2xPtBCRl9QfPAnT34xMUpzMfvDqx2QEgeBhRXjhNm9XcRKvxygU6jGS15Q1k3cBpYqgpdha4J4
NTwSUCIqLCUAofMrWc1IUxzsgh7UY+y15dW5FHhp9vJlu/c/okCv4dncZq2WxAHvCjqaK7n2R84Q
+y7vkp0UvNiduMA2hFnVXFH45WNu/XDNmfKFcWzUnP0vS4fgkPUfezotGrYAXbro0eRDZi0G7bPn
7aMJ4UiETulHFaM8dWEg6z96P5ClOwuzcPd4czHffV1+eB+K8acyfFcKV5WFdb5oIqAhHyOs3jDA
sJRg0ibnaPY4uPrAdfn6eULVl6C3S4N2OGDx6yu67IUqtTx/M3Z5h0YYF6lJFOEtcABtp4JytwNt
y9qq7wHEt6GQY4kPDHl4Hcq35FOQIDa1uzosEB6h7/fk0ZhUixoqbvv81TVy4vXiHcXou894hJMW
5Zm5NfbnBjRwDa1XUhN/AK+7gER4PP4VHT4BOBwlfekkF3ylvrZVb1nzUFFJnFmLVBu1AcIv/+za
Cl/MzUxqzXZkDgPAQjr0hjDa07iztr7z6cZgfaybQs3Jkk5AIwe1oeFeVYo58hkbR7umzqOPd5+z
TxpB2fQhwgxIz+djkJFd3MVtvaR/dNbJFFaJ1IHDQHotA7XnSepY0WLyRmlVOaLSfHfNlDeHPy+O
5q3b5auxFpaoM03BVZ1TiN1KAX2wUKf/SBrYVjVycGYxMxKgq9Xk6v8CKa5m9NDUQ1eskoj9W5bY
L2St8t0v6PmeY5G6ocud6AZDI/8+stOqXAbB3USLUVMsz0yjeMc3sj5Qbkgdqi+4uYmh7G5txIeL
q/O8BWL44//lRlPwk0FhX1NiWhXlllIaZtr7XxRre1ALFcUKLlac/RaNQvf07kZkf/aut4Gg0TEH
77vICFwGqKRwKZlaRo8tzaNRyX0lWxvg7tVWWwkrMvE3oTcGKKI8RqnBwatypK3S+AWIdJPa0ppi
W6cdHzDiaey8hh8x3KYuKQhbGJqGw7JdG6ClD85KA5vveK2vHuLlQE+wEn2NpL8LlpJvJZ0W3za1
fCzA0/93IigI+JEcjKwu1m8+R8oXcgqwa6GeybkYitUK9r9MEi9MGDXAyEd6RSyAMwSAekSBRKyO
9oqprNrr2py6mFzJhsYovHfhHFces/4H5nELmrRGBE1Kdh2D25MVfn+x1Hx+i4XmFHLTUdd5l1og
i8DRxeS1NH7C1C6U6lN2k7kyo4WuUlGpgCVWE3AJize0UjSrkr7qg3OqhWQ8uqB223GveDTe+FBf
k+8bwmO3/RRhwx5u3v0d1MuunVu3jw3dEg4x0rN36x217x2jtq3pvJGatnIXTYzR5KcLE9+1oQKh
bxIVzCeeDoglcMpHtBm06PWdkBKYH2biky66bzTv91+3uPL5IXha7HWhPwkAmFnyM9akj3pgLTmv
Odx9iyS5dYQKMF0JY7x4wDxv+CBJW3E2BWe6ru8X5VQEXboAj8P8onCmWNR+m8OOq3J5s10eYofa
8RyGXSX7Qc2um1ey0o5mbRwIazjsILVR6LYPV7Ry8H4drB07ek97Qcm6N1ESx1l4x0UW26FMZ/7+
JXEdUy/qsUKsPeUo1bLzte/7OUInNIC+ZlSHcQ44qg7zkAd2y4B1ywd+G960+nm0ZvlWc5t7o80S
tbAcPdhdbnUjb9CN1jsPswlOtxZpCQTcU3gr29IaRWid0tRR/NqNflEwQMB8rtoA1nsgc9S2Fulx
UHXsaGFmy31QjQxeO4M1pPIkmtDvzpMogg7v0CeU2rWzJOqd90JwVuLGfYlXsEv/4tEXgkUVSOgX
gRvEqc5hRcB0SAf/oFmuN8OxfYSwdlJFXumeM4u4nKYlMb8vj6QmvxaqxqGNe9LARrC6167ExqeH
mgovP5Dy3WGQ6fg405Tu984ijO7kP8UM/tF04cogUopx6L5dC7f9BEcPK+W57IneCO4FpzVrHJUV
4ryNTwfqPRy+BS31CYv86itpYxqbTdxA6av37pzmeomYR6hoM/HdNEtn+92bQIUP6oBzbWKW16d6
BNFeJD5L7BhXNXkYUFX80+89S6apZxSTacRt0Ka688Uc5MnE0GmVASix6rOthLmvZndIqO/Jb14Y
IQZe1P+vngcfOa6R/cZDhjipv58tVzzSzJTRgTyuNB8BT6U45o16q2ZUHUMU44tN5+fGECc+/LW7
63u/8p6LRQOMYCzjKsFkcmCA2rMvrPb6E2ffL07Ofu4vj9e/rNOkOqgVqVQKMI7+FESU6j5ZoVv2
A63mJOMJwi1MOaids07KGQZxN1bEhSN1bH3w5vyS3c+sk6rdKLzfARb0VlZjA3LEVZ8aHV2O+x9r
n6rOj7fIHLjQl/CMBsWP2XBrzpoolOEh3uzG3QcOJo3YjEBk1bIH2ipaCFovKiIe42SGzGW910Vx
9QG1B8jtQY+IoqDzwBfKDyJhxzxiLeET7Pfhpuwap9tNsKDuZcJEtq9kcYFTgY15m2xx08vHE6BR
DUlcFr414poRiLeU0A3XIjocXNWf4S7ag65GI3N819PU2Ilhsaa/wXRmFfbdWvl8+MC8JfLe3ZbL
ukRfVO6whSO0Oy+QicN0iCD297QGyrLnCXLblpZifFA2+qmpctsiGHX8gYg1E0wz8tI5iAnjhZxf
HY4n/SsUsM6P0bv7/Hj7m4qk3n0enVW18qBGU3C4U+GF6v5ilj+Rrs9OtUurAHJibBw1DZlomMYF
+conYFFluYXAAHo8QtqGT7pEaYvmBJsiRAeFBaBSq3Oo3H1gNhrOEm2KaAV3Xu/oh+ANjix6X0v4
iaVrFe+YgZegbU2dgITMvvx9IpxMkowRYv8zCRVpeKOlVwjGUMgWJlNX5aVAwqTAEVP2YSzCmR6c
xV1Dlmts0H38HbgtjZM/DA8IKksjg/9/xikZxDv+dqHCCxV/MjSHJdx2ob+t6YGOsEoz+ytP9yEX
972j6g990X5PdKIdxc5EBVHu5gu31CtS0L4nQ0/T8FMzqV01ApOWj6Lqy9zcxf+jvidkZJGUmzbA
P/HIFQmDV16Wl9lpJJz86X0aqBuLrJu0ZVlFfWFCMeM3MnSBvaWw8BLVlbWTtrnGb/T0MRfw+iBi
hOLx1+L1ccz5r55YCU/Xaz4B7ZFLGPAXKIZFh+VcnVO8TZ0A4fAu8qD2EBrjn/+QtnT6yjobonOQ
Cq/sUM4oOPZnV3hTM/cUS/+LY0Yc2GKU+K9Yl+FY0c2CO8FjptzNytcavVKgZnNB0mY51YjrpVX7
579k6TgkpAsxFPO4QfkLWfrLroolo7Ri8K8tYsepaR4JAAXRtjBH7qlWtV5TNqMipyHMjkdkeG0Y
HdjOZaT6HFoespYU8EGdWV0bcf2eQDvj+fOnOdieUD83H01gVZ+1eD1DggoNs7kbi5byyXiCPDqt
HHKiTfh7EA09A4Wpum6/gz8zOoWVjobcsTCebWWgt1969EFLSOmoEG5ISGtYEiuNGDbRbrwF6vAu
vurwyNfUWnZo+JShyLW2RLG6oD0WsPNlOeUvouEHvb0mLr8kp6zs4UBOPHJ9cCWWlDRKjNNdigbS
EXvsRFZGmub5M03YTeeVu6Cgo9xf9tFg7LN9sCGvh5KwGPD4we4Ad7+z5BqsuOTK4N4yO9q+mMKi
9y8gCnTi7Z8HYNkytDpWdmDT98KZMDfsv6IgcwWV/2NxOZ24cVl5mO98NtjQ9KrMhXvoZckToiXr
JNOaXyQnWhOxtLbAQRGlxf+8RvnAbBQCaoKxHiXLAt8BGisbpyGyNagzGV630Bh/8ugg+RvxvTdT
e6ULU2FipY+uHNSiLUFr8hOKAxJcq5smXWFwGWuhDIvYSnMElRGLtZNdXN+x/eg2+2noKtsDLRnR
ytlUNakGiSO2FqJa497OIoIADaU60ZbqzfAOXAfWHS2jwhv1zOpeeg5HgcBFZYnqreAHGGxEzaKk
Gys+DSb/tWuqOC4y6uvOOkiflQLf1OXZL+f3CR6iOlW/qZJFTSQFGBIzP3r4MQbztsC/G412Pt23
oh2C5TJM6RoLte581na/dZiF6c91CTrAGGdPjX6Yl3UMdXxsSbk76AIT0+ArxjDTJU48STYjiIoo
nKhu9t5CouwIPJr/qESuVEKDHFFshDRh19iqdhndvTl34dRVADy/UCpDSsCk6pAMYV35glk7eV/I
3CyjDaFW3a5bOwxrkeIpfgfaPKO/dDSdKfEmfUca+PSsanV3aXALCvLmWYCucTTBrH2Hcel1CJdf
z3RlP2RGfj/Xv6TjYE5XdVNDq5EFDU/hEZqAeyt13wXnNjb8szaVs8B8UaytNB3sea3/RuU0jOoh
JYorcEXpUBMPYoBjRULwoniU9Y6V9S83FSe0n82yqBow6VaLGdsSkZNh0fNLitj9mE33lMFQEsBZ
Bda5HjJ5TSdYlrglygpiESuWpd8K7cOq2lrKF1ElPJvBN2hu+1R7cBAgXA1c5tZzn5ssVNmzyXu/
upeFgBzc12jx9mDUN6hh1AsWKRfo3p8tUp206T7UwPVwjKSt/GK7rKe2H4slhPr4FtRXiHYG+G87
uyHbIJ9366gpspYsvo8xK+pO5nC0FafYSKZMBlZMULY5QtNEMF8bJodkyoedHARgma63iR+nCRsM
qiU1Ewo0ldWr/2SJeVSifuH16SrUXYSm3bskrp3pVZ67pKkut00hCnWpGJ5EHSbDM4Q3qAdyxhkt
dmYtCWAbNHRwDcR+rdoU8rt/HqhhaZSsC6NUzyGpi8Vb7d+2j0R62m6zzkMQrSBUdD2biLHus3F5
VQo7i6tJq7VRp/p+AbuPFLosGSZBXxG9cnfYsesejWOHOZF0Nr9AbF/qtIYtDtTYmc5yP1gRlEPh
n9TXt/Z298ADA3dWRNqVWpRuoyiXIuOkaIpj6HUIZqVWlHEOuTtH2cj7Ru1NFtN5BPu25oZLvEAK
XAhbuinvtB4Ibl2Z10qwQkuZ+/hQdFON/IO6oslu+whGD8/5xp2rO1gGZTd5b004N54/yhcnMSkF
eKi/HsRrjX8WBrLmf4qXggGeRIwCYUBmu7IeIg1N3wdVNvhZJ/5rA+Qjv7IPBPzSOQ/XOPS+ULZ0
Pa2iV5yjwO/U1BlmTF3jeN3LpNZQYH6dGC7805fbj5YdP9ckwfKp0MoWWOfMB0FoHf1tda6cSjRy
rEQdDjdfzMV2rwbdxeEMZgA/SwR/V+RcDstuxTp76ZzJTMkyDtcmtdyPoC9XDUqUKGxjDuXrR8Rv
YvWyBRPW/ChT/VjKJe+45vK8oiokj8FqB67CrxgUgnd1YCeD345/ResxB5MmtXyPW1NlVmMdZQpC
AJlgpQdO3PybVV3ObU6Yl3Dhb590FaVIvHumzsZRoNnjirkIXh2si62Ny5YOpuydnhPr3GHPhxuN
yXVJspMyvyXfE0ZLLi8k3cTWpgZYOcMTz1P77QA3EY6cFlzyRGgQ2cJA8kgf4W1pAObzaJ7o+D2M
MESo3HhmFaMaQJRB3AEYwiUeOoWPX0sr95juk/OSuen0PfQY97Rz9VlLIgjTce0XrU+n0bHrSf2X
OcVwcHTb6Q+dTJjtgHdhKa7DwRAdCar6EGopPYtkowrUXc8aRhLZsPknHS/oz3YZ+dHlSslqhshp
i3ozQD/aWX9fQz3tJzTxtkwZvrashSqxt9JQbWle5Gri5DYX1fs319/3M/lqI00fekwsLWR9DUWt
Xo71CeJ+5Hzd5xzuROlx33zotP1jesFGwK3rtdMOCgZdiNg383UHMgHi4I5Bav50Eijs0Wtq/IpM
k/TEArh/Qkxw+fjlglaMCUzLOJnPGe8yEQ7K0VWWvLQnAEnkDqs5hGgCuDESaruah9ch4BLXRw9u
bHQF26hPLDRP76b5J2nVze9TcURHNgK87b8scaXMvRCiKne3qy4cTbt9CfPocK3+rVDOAf8bBlYL
XmrE9wrRb/Y1cx5ADSwZZ2X8Jub1jNskf72OvW5FtjsNR7A+dsnXlQ06wXb1F+tbXdbVkFbxs9MZ
d4ZmBeR5dPzljhcV0Fy5X8nPGmyOMmovIYqoRUPdROju5yc7lWGL5stsa6OAHmnM7//0DR635DEr
kSAcr/+nN4lIKW71BnXPwvrFrtF6A7qFrIv6m0tBbjHvmXo2Aljr6SrHx2/MZnpgI/dkzZK4P9VC
bkOv3nmM9ESC1DRpIS82yDlLjouysAkOmtJYs3W/1rDm+FcxckoQjMFTX+F67DA271dwd4wWUz70
TTedINgM7m5wKwbyE8g0oHuakGVpnj5LzMolcgCXhawR8T8CDdnt2pfOf46usTCFI775hBWW8Vwv
K63He/C2Dzjroqb9IPwDQhopfPhNlKJcrVPjtl7o5ASOj7Gx/O1B7BKEsj5dst1ZI+Sb4+jpSc04
JpSBYYXOmZx5uVFemdjR5X6IeB0UTWYLdQ+LsAOGu9IKRaxdJ8oc8l9GPgVtgXWM+Uq8OnJKcomy
zSuicvIXYD9r3ovHd19lnNC6OPUF4MTE1WWgDnSJD2Q2jN2nS8SNE/E6NaXXVqyv+1JdtKy4ahZc
aYpVr09Vels3IJZ2YVmJpNoRUhiK39T+5jKc/LhJLwlgIV+6DjCC8ZqnbwLBUMvBMqDWvXV6Ei80
Zfu2ASgBsako3UJHPPjHjnfGCrNlTS/EITryghQuY3qUCAt0xK8TwGFLTzAVOTUhCmFxRNUr3KeK
UKFDhw8m/4cYHBlfoNYNyZ37L5Cd2f4YbeglScUumnfKaemPhNOYj59w+lUnD93CAPbv8D8EtArS
xB73fZH76uejqpD3KUyfnawLJ7nbUI1WJOjPS5+V5XiDWAKKJL1vFctPhIw2RuCpY283VrgpGFXD
Uv9FKRF2y3++0L7brxESmov993eUZhjbv42+MqFrMSk2G6oDnH2Q2PpLmFkGJ0lpNHxwkluMlWbC
Kk28CNEnQsTHMkMlxo6LanvKdnXVjuiiJPnfq30GLFS409g0sUf7X18ZlLLxgoGdkTVX9XSxW/c5
Lv9cxwSJ0hLaIvxoRjoKo66pMWPBd5Ug9y8bgnVaOgJ2Qz64FvaoAVnGzvJS0sCvh48ubvONFOwO
9IE4BLA2PHlfpfGvOBGE6AlaGWQwIDXKFLyqMbZacf/4xmk0xF3urhZmk1v0EUARertaU9IfzNgn
42kKFDAuhNresjpwWZK5StFuNowMcgoLEN++RHRw6A0gDn2HxD0P4h69RlnDuM3girq/huyndUYN
N6ocmk21EybNhkZ4ZBBoyR9+GKSsx1ZRdQV9unJMKc9tnrQch4aHkA5Nn7PBqh/xhUfPH9XEaCZG
1/agsjxbf3EsxtU0b2Dli2PbQi3bcKXToQDj+tl7Ki7eckE5APVfDAVy/BUxxLMOj+aLWIOjxfD8
0ud0lQev5081MOHDIoSH9n4yq9c7+bn0CK17Tfq2TmIFHtizNKrHdhl2N3lJP2slnBIDJjj8gFKU
vetkJQee5JZ+sdKVtRDinrr6S7aZIV/hS3N5Eu0Vy2zbbUGozteHPF0+E5Wc71GWGub7G166DTae
8OVeH95ygRj0UUfDwiPBkFXR6DMuhReSbFP4mkrhUBy/QjNFYXfLhEz4pn8lNt5/x+vrSJgBdZ3+
LmHHxHnXq/COP3nVC7Mc+OaA1WRM7djy6Sbzqj7tTHSwEEH9YktTBl665cRWGjV17YKjk+oBl2n9
5+pmgGf4QHQrSfQUbAtnHSOt7v5SbpZ6Ewkc04Q9aTYw31emvSbRDRvaSAdi/bXEaicUc7lenIp4
hWf2Du6i2kv6NBGDCxESYUaomOXpt0WGCUMWUCgm3dVMGOCwGUNbHgj+jdiQ4X7hOvaY55Duh278
gVaCGFHSEPeOMS9rUZZixDpvy7ylMHHPUXY0sfb0ug1XiUg3oalruU/NZADXDevyuqtdNyhVvSxk
a2SoL9ahoB3JeACctP9gFvLX26wRcgBZ0bQ3dsWU1oaUfQuz3JpMpUsenRLUgTo2hHWG3APVf83N
GWJKSBKia+oHXq1l3GdI4t55wcKcIcnDTICo2LNx0t4dLTeZuWSfU55gfc2HJti8pelDmd2uCxne
a8tFpfcU4y65ST8l3NHZQn/NPj1iBSsYZXBecSZ+evbD8B0wi2/wGtOm1GBPTFPtJpprwEK6MOkQ
tULfWa8N8USG66RMkGl23RU1lZ8Z6g94+fqSB4tb6Qrr4mm9jcMNq5zsmvNqoijA6MJ0XcjK5Rrd
0zyofZrAq3ZP1lhzn9NZble3ppZrjIyZE7D7/BbfbEXJCvBR8Lk0c4ftQDzY5fpTOiFmZ0mPVWzJ
2htfNSdgAa/JZsChSrtbGVgNmxH1oKW0z2M5oCAB7azK3o9pObV4iehQrQN72M60ZrV/ZRcrOkAC
ZmTqcge94ETSV1pBWql4DNgLFBcUTKWj/0XnWigtthdqjZmxI+64bBVKpGce/45DLblccPCpzjsG
b6Ljkcmil/RTlUhInwAJ3frOcY6reQ4l6gIH5ybOY5zO4VxbuWIMgB55FAGJXsYCCBS/o0S9xTgp
aJdF7TSke6SyDC+zzytMXNEbun/+cKhuLI0NQxSFPBKLw0fAVfkwxIu9SElpS+dEu8L7RNy01UN8
vw1pGx7K3PL8BSgNbcooGp2uYc4vEXC0vb2vcL/1zRRqHjJKHSe+pammUKBbqej3JZolrJ9anBfy
/DH3FTim9I4SrE16gYmeRam0pE9r5a4DhtTfeoAZzclc0aLdNSaFEM4k6D5BMJ2pFKp1XgAnrBgb
UrckYJq5xfWSPnpF0xOUwsVFkvkYDzuJdPN8dIeLTkXqUfAYPm2Q8RftL1tDbAqZg+lD+DtkKRwk
35Wz8uCP2jELA9dpvs6ougtOGZL3j/eDwsEo/sCV0CmiJyO66Pz0+3Mpkt+OeEGm/79OQrO82hyj
/W17Wr89oTYtqhB8EUQN8EbHDo50TORZAFWD1GZdyQYtp6/UHoVR5LmQRN33hB6LzOfrQ87zU/F2
P/qIQSPYQEp6UjP4HyLzXAaxhyaoPOpEMSCl4lW97zFkyxMo01mMEE7Ow+fHANFWX/fHWv1F//Fb
ibA6wvg9Sp4Mc4xtwdSqg97MFvIJSKuvReLeL24zsd8GvZvPdtFPlTi7rQ7ipjtBf2oqhGNujXo9
YWlgoRqAIkzZeiqr0n0eemic0WGhTJBDN4M+s3JbC1FjahsOCOONrYJ1QKhK7Xl4r2oIR9t6HuOY
EPbpmoF/Nhkb9pQI94VSyODuaAMPU0qL3uiVUWIXhLCBvdd7VH8BqsAEPF7IxlYzwRYCVEvpy1k6
La2Q20Zb0B19LKi9TGdgNiVk8jzFcLHFmIT2tKwfgOXaSL5/F9pMD7X8QlmzwY3s2inEi4x5e71q
Fk+WJar/huRt8xaT9nqqRK5+KUmKOVhupc/Q7jiN29WZ5RRL9lAPto9ZWHL6kBojbgeyw4eRdk8T
yerAirFgHeudpmGSgqlo6BWTepEGXG9fmVdpuTkxc2x6C0K2d0rw9gXwWBPawyYo15Zw+p2r8E+Q
ztp4OsCcJQbOdYi/ZU7HEd8y1zYXH06XfuhkGGas6NN8RpQT5sa/h3Zhc5puk18+ZKoGVhVfcUHP
JZLQhlCEObrD+h4F79G9QIWuETKI5IJxEXCmgg80pIPR5ybeO2t1HuWEJcbJe9rvSIVgXK094sip
viXsjmkIp/+MIf6FHftmTULReqAMC/+qoO19tF5/cOKbumRE+1Ne5WbKYhpvBb7+Nhf3BP2ozDCa
Dl8FZa9v9pDk/vEB/AfQILp26JFu4hexMUGflzfZqECB13NQVyV7M+lA+LbkiKt3Vpckc6SlW7qG
WSvhK+AhKvL3L7rI9s6j0VVOMuq6k5g+YJP5asKArgLC9bqvyRZ1c1gb0i0GLJrvSIescWYeisBm
nAYz407ltTr+LqXNhdaMv3b8h2JHC2WNWm6MKpT8fNYfZqT2sN5Cq2pfnaEyoioBzy4TWRyEP2t+
tVvyBhe5tlnVmdKVgSjieKhUL/dB5aXGJHdkodEt/m3sgKJk1IVg9KeGweHtLJYJ/ndQ18Nv1AoK
DTJlIfkEkXkGtxlwFGCMpLjw9OkuvjEjA/iLWngudJ7aPGDQuABdNw08y7e4mO7c5w++ph/CQ8Mp
kTw9UXALXyiOZz+n5ANwcJUISaiWtw18ZkAIt0ywFi7es82YoeYOoaIG8il7uQgMJCJYu3xFVCKC
yCqZWxgwhzA2OJrtwIvQHJgN9AXG2O9sbxs+I8AL4Bo6dSm3nPKJqF3WwrPenGAo57sYpKAcK9v9
O2PQPJMQZP2GF5URzfI5thiSPyDxtogISTLZ2SU66zP3bunUszbD7p12ii/O3LkJNO3tNwfmbGHK
yjpWmYzoZk4ofvsB4z7IRLkPJLaPJ3tiP/QRDN9ShM0kSkvJT6Fmw2qQyJUIMbOdHTDQOit4RQw0
KqB1GNunH6F+3mRjw449msbJl/C5wb0zh77+OQJjVVqDjF2iWJK4wYMr+oYSJ58ZAG7pF2ieQVCY
ciHzH8nXz0ldfyNoupbUwwV67pHtpdsuHe3nIvKGARB3UF91Aw+KHFmv3XwJ/yg86WNeuiSYIwsy
ZOMGUsxBTqBHK9yhdNEntWYhYu6Q12N4bSH7C32Oizq+ZGG4W1GtcNab+R56D2lqh9yfIImdYcyi
Kj9DFAYShLyFd9GCcnlOziGJGBkdteyRJeHa9ZjM7fJRn3+oMTzWIMDXfp5fWLZlBc34zk6T3u1A
bgwaxEcjnchul6KBzBJQ/7HpzCcPaJ8jRvlI4PuKI+pIsY1gnVowo243IvGD8wosIKIHM8XoqPHd
oNpxx22xM/eO793NbpBPepEHYKbEan8JE1Ddmyw6kmZZ8y2rsEow4vNKWZdUXiKC5lb2hLtOAgIj
Hjp+xq2/B8RBZx665HaJNfZXkTTs0IyXpJqsbWASpFbwMMJZH0SqpKoEaXKW3dLMUuiSo7Ol39Bu
D/xsFUqUdYPGNqD7gGCoR4t1oU5ejbrgHBsxCVqbrVztpCD6j5WhvW6xYopTNU0SZHNicVGgCNkI
Ti4zUAwkccpOWwKdRNfkX7wQy/Ov9b2dW+5m54CLV7+ongGRph4byme7z+Mttx38Fs/OnHR3FtqI
LqL0lDbwUsJLqhZngq49ybe39SMsnV8CN3gXaEar4Mo9DOmTjJQ+XXjyWQuoZ4Jo8A3oJvztRQA6
yHggYwVAjxJpnlr5/Aq79XrCQjYaJRL4g/KHOaRkES438/1W3MKADQDY773+1TGSVPgo/D4CYyf3
U6rA1+nxTLdiVDy6nLJgrIHOKYDfN32Vmea7b9ayHtNXrn4gmyPEfF7+e5N3/6jm/WZHVeo3kFeK
hkQCet99/ekxwLu+1pSOqAHs38BH93pM5NxOUQz0t3KxrBn4HjutyIMsW7A10t2LJYZ3fnLEWVpP
7Lrw3NPkxSHzFuyCtSlRqDD77Yy17Tpjlh1uZX0h+hzzLDXKh8CHElx7QhioebZxUy3zp+t3f/yv
6B8jWtuEGZ7492eqjUB6ptR0eHt6I/rp1PoSSaS47CXTyC8e1ldxlZNUtsdlbA0OhrnJd76mm4Eb
+kJG9kNxvrdURLGEjivlvO0259q7lkSdkxyLUoDCjgn2sHS7Z1Dpn7scRKC6goKqL9U0eqXOtM6X
efEkSnRyosFSLSZdaizvVhvtdLwlSN4RKzmvqMnri3R2g3aiolmQBCYH3/Rigo3J0MuEWLTwms+t
4rnMhoYKDVxZu0Zm3C6wJctAlYXzid0StPQFuMS86AgIX29x2dxF1YWpHq3V7OT+lI/FknUJpV8P
QP6VowJ6194cGv5a5AT8MAeD10ApEUS54oH9Daxb9PnQzHYdEaO5J2oQF7tEyTHC0XzJukiUgquF
/r/bVEvKnrX8/p/w6FnvbxjC3MXnjZzwM0Nqgm5AagiiJBTsOhE8e4dtuBI+zZ94BpHNTiDAOvbg
fgtitTLF9aYpEIXpir4JshrpWX9/nF4JAUxy05TjAIgxhqLott98zTKUsOR8ZzfzdrDrKGNdWkF3
2hC3dNqsBpSy8jvVS5ST53FvI81pfWBmKFJyoC2uUfuX3RgpAqR2MsXU5zkd83KQhYJlTSO4fmSO
qymZ3OvRfXc6VHLGFGA6Dncf2/YisTBFXIzhx8NV/iiPe8iRS/k/5CdK630/Pq7DQTvfiLTZu83M
ybg7+gbHmPj0pUfjrD2XJDBxXzZRxUzx/vBn8PZeBv8MkhNC1qa4yrreYlzvGDU+mr7dgq+1sPu4
afikyCZaz7OWaShS/REKpLEX5oPmI4Ja964theCjg0t2ejzs98gZTzbBBxnRDYpZGY7ULX/ZQQFT
0zAFnIQn8/Xfhu5Cf2y9SAxznamlIZvPeYuvb7BHYx97IZUBoUB5BXsvN0eaLtuvLiHKR4zEPARO
a+pfCx/Pfml6n8tWZtEg+kWdAa3PqZFStzzFf5lk1iMAhWLOJ6sHt4mSNlJI1ObApy2Rs/pQHdGf
vEqNN5Om9+Fq3Ph+ansYe3gUXk8OEa42WLGvzMF1rTUXtyz7gv0Cmf/dYNQGH+b4AtK5V9l9OUwo
Lm3+XesGjvI7+R99rWXGznwD9OOSATYX85KIgx2NCQ+UJqYfosacARt/VhUk774mODH18NVerGe9
MGRRO0KcV7o8yaqQmQfp0jiaD53aaZ8lqf8847faqVeEuuGK8EKYhwQXPIyrdz/Ij3ou5o0S446p
Dm5mS7we7ndEJ2qL6RszODQFk96bqCLfNKI8jclsAD5T/GHFCUkbqR0r28Edieb4jnNh9J76MdJo
uKijBr6dkwBflbJF7Llv09+52Ay4cfOvL1tjtJ0ZH5lnYXgPPFApJTBOnO16KaYy2gQ+qEvum75F
KquFMqCktHuAHt/HP6IoAQRB7uKcVWkZpFaDZ1gOtPlzH/qhZMFOKwvymNDthO2LrfCTXoL49bLC
Il2uSE44/4jXctbmS+r4p8BmXJdoEAJ+X8JDENzHQ4jdGBag8eauazGPj2K3mi9mmtxGankBoupK
ZyJMaEZ+C4UxCCyjaY7YaYSGm+VHBMsYgcGIBydnMDLeZa14X1IyU/OH0/BM8aGf9xIfG8O1/MFv
N/jW9qp0XdKZ/yNk2BS3xn1X+0/kAT60zAltqmX36WDnLcXMF19URH78hopPRRmc7YTbUlILSTIo
6hQbyr0LZGJyYK5+yznc4z9TEJREANq9DGK33Bh8z/8ryJTUexLcjB5HtYVQ6WAoNhleiMDfUgXg
kJak9xOE3bHI7I4ny8y6FnfLygeFyZFqE5DgaTRLT2NCFWJ0RzDtqTitJd5g4j5CR+Gl6+m7lJzI
tO5paB9oDfveTIvuH4dz4bufVxZKTy6t0STp7JsuTW66Nhx4njTX4tcfyCJ7ZgftzoqxGW502hY2
kv5G6Xr6FM+LdKbY+vt6U2nEZoVJmsloK2xSX1KxaUbStKiuxNC4JqX1nXMYbFTiBdAv/XrsbuOG
3BzK22hO785b314CqcUXe18cCw4BB//uckz8x0H1OTAA9YQAkIAgatyC5gtLSvaE4gLnxH+g5xnO
zy++HwMcC6QLWWr0P8mcaE7WK0B9XbB9xT7jkU4FSW8G1vLRnQG9dLGpXveP9BSD3+AFDVOylJuT
L9XRu7zyAntvTeGrgrIUwaqDFcumu6mWE/nSp6ObgbsffoPeAjWVA7Qhytss6Cs508t4wl6oh+L9
xNJCAS5kDiLn+HuxeEjtO3uVy3jtnh4SKXbfr4ObZnMYTPD8D8EjeVoFvWWWtOtmvKRO/yh/Wk7U
1yx0bc2JoSVLDoRf2dQp2qSdPizbun0z2Nhki2gftTz29NlKdfeaVYLf0ya620YENI/3JI5DHG5m
mwYtSyIRY0PH1iyi6CVyz8cuctRtyKLex7xQQ1AhgoLFWLGS4Kw3b8u4CYsGiyQeY/BXQIoeX3cp
nTS7qDKau2Z40JtvXys1Uu0tWikykbBY/4431evZuErK6vEO7nuI/qpkXIWGPw044jd0F4SAc0Mx
ZCYvzP4laFHpIDm9s8LGNZw1UDRs0hrOYP07iYeCOCg31ithACzmKzqvy+GbV6ctuBC1B3h3YpEH
gva8A/SdlhwFps0vT3IkQJuu2iH78ufLRcKo2VrZDU1MHIEsatha0Imdzyp2VM8pOpY92UqFUQ7m
/WevBqlEd/mUOhy+G3InUyvpgXNIOyXeyyGxBzJvsXDMU/1Dijwo3X8nK4k+oklD5PPra1/leTcr
c43Sn5RjypMPnRC4Ve0v7ghsqiNGu3THcZ/bcEKvuT0aT7wME0KFCJppXvy8aGD+AbiD6JrXRHDN
Am4HyS3aaX0lj14CiZ3MGIZfiqeHn5VF4GOyY3al+BFiWdnFyFDQr0UAD/1VxPnTCpTcvw2cxAOu
OMcEluP91OvJIA5dTGZvtKgins80Qlp9zdzAEPIZIOSrwCY1DdRfum/PF31rj70fXkKCndt5Koxi
abuC0aVRTJe4Sl7GUlHTpqfybMsofTr3EktHxsemATImPaq1vJlN4enyOTbU5FJoNcnHg+SvvQrB
+L6i1qpAjib/OwR8O0Ra1SjsgYLiFaHHe9SPLy32hZzncIuIER7clxc516SGY19ig34TGp+v71Kg
UZ/nzk3ycSlGxiCbNtKiJKa3Aw80t9XBbEYTEhLaRA9iaPiHO1x444uZQJ6Z1gkk2/5ge8AZIwrW
Fjy8HUUIpANlfutjNzVCvDInmcZ4sb8URbzsYUfDPIDMHSoKXzfyOAkBjZCUmvsGznXbHpTET5E3
MsuqHlbakbtDd56286cDXXDRkdfVCAqEbl3TwRgGfXBjADu51tFzcK4bKZ4NPOiVk95zCtJ3LLZU
Jrn6cYh6sU+l2cWV3SFv9wqOHUFXZQt0GH2nhMAOY46ZyUtFi6LcKxDgXSgwt+3gGEFUhM8AwzGm
0Deg5nWlbVAb9g7jj2ZyAoD8h79GWS2nnpyC3EuQ7PO+Y9+adorqjcokMnBJ93cnrf6otQC3jOc5
1aTfYydKiQ4LEP9RvQZJyE44CidWxQzp9mZW/jTaf13auEWZE4aoVlTGALwq7sF6wzwgHqXOqvcN
ed44yZYR9pCGw3LObXoESVvSqubineAz7rtpvx+X6/LjpkhGlFfiN/jFMypRh6nSL8uWi4MDzXYz
M5ThOfGbGcvbVUJgoBeG3PiL8OH0oKyoM0bbQ3gXdAqqJNAAWB7TPm10hOISqpcau4TsmFf5Mlx5
CYf1JHLa5l/X3MIW45moFZUrRaSBtMCw8oRTaum/+fkMo8z31riOIMdCD4qiyqTiMo4+flTUYAum
lB69af5YeXNOQ8N85jen1vXeMAjmaCOGcjI1voZI+2St8QnjheMa9As/0rafNqTz/ZPcSOMa3qMl
2SGgE3frMcYB8iN6VSgdIidoBjJxX33OOjfWLP3nNXz8JSQz7jOr3ZHBFYb7YXhqnmx1iZEtWX2G
UkbbG1sv0JVKkqlb7t+5u70CkZbBRiKPAugEBo8622oYucdKO3IiQJdrwsOLFN+bvReaqQz3YpDA
wJ4UO5zIrzevpZkLkRvonPHA1BFoAyczQgBfSkFpDHzCbw4B8kYUvV6Aj3K7HHhmRJcknT8VPN0t
uE7omlb2YooufG9qYH4qiWf+Y4aJ1/GQbq0nNYdiKFCS2pRQ+SWY5A0k7b5ILMdgOb73qzwa0F64
PM+1A+YI0BuirBdYXsHtSn1z7U9vvN1cgO6M5+RQC+w2GfAMw7gJ53iVJ36cEXyWSfBP3kNkZrHh
BXdyqEx/TwDidwP2KY23a4p4OHSr2P+daqcp7m+QUmIF5rIzOU7jxqmRvJbHi8IiQerNsoOAU5Wn
xJ0Dd2n/J+0ze2/EeCBGCvchIe01tb9TliEqN7TA8F5z9AJ6oy1V/IYtMs56N6uUrO9GydNcDjpd
Lobi0iQqb1sBbRYO1AgU23BJ90JknfMY/W0/zmXUyhhLXubIclH2AxO2C0LhgOR5WS5dk7Tux4uO
js4dVnYEKLUrFs2+qns9i/Gq1hV/159ovaNBBiK1bIz6OuOijhYS0VcMKaHCwBXtOGAGA80mbjN0
bM6OXHSJvKweHd/uqxsGS8L/W0FhXBWsF8+L2NzTVdSyWm+A2Hkl6O2txtBXPDF1dFh5gSHs2Zl1
2Bl11Z+hNXd/Ozrt9AubzaxfMAiOfpqDeIu1fms852F6tQ+PAc12I6/2YqbVoBGYjVz7rbiMSShL
N5OKFQSTlq24ngPTKchAHnRMVAVpiwg3DOrmcgXSMZb3+732X64DO/2NGQ70Yqit6/pWdg8WDPeU
xBKoVLe7TRos4B5PwU1O85/2DJTfE3oDTN5RNELPnXk68pjwGML/vxAc1SPjrflR8cigJsLDpCHA
M1zufZxkWF+bUZU7zTa1g6Pbp3AtCAGQc+Tr6c08rRTuNjBdzhVTiBkzGLUxFu4yPIo6tRQkSD0G
d8Xlc1RZ/STHw5d4cS6wRnzdDF/WaWOVUMtKkNcC2vpDAX91ecj3RZs+jLBgMlwzs82OOhG60Vit
T/HvXigXJSNZk97fjcP1M1pGY+NTpZGX9P/Z6Y/SCYjozDRxcxdKg51LOlMtTtueFMG5fdKKG74Q
FKFjjxRi+3NT99vcrdvY1xqiiCQLR0sU/2UNNxnn69uq3SCN+WvtifRU3j1S4CvdbcJHUOshnJSv
U1JrDE2IcEjGL85QdYosnGqT/feI1fdSdjSJJ6a71Fyto2qvYJ2WiNu6nmBfZ5IbOtMEJHS1GRE/
pOE8hS9wJqHz1Dy+aniiBl6e2GqHWs0Nb9/sJAPh50LxcQTQYWxmRBI6NhVpdYO+afqPgjNPItky
IIb1W3iFyNsFP/i2z090/DVFXo0nsEqmvXFSO+Izhv4BHGcFTVcKTAWTFzd15A9qNeNIqcxFS04j
VNyWOjZlRrCAoeAYCTUDht4bEQu57Y1h6enFu2NF+nj2gicJEf0kRR/kpyw5zJQj5a4Mk1JBMBls
X4/9AGC9oViE7vWhaznHR5Q42W3Q1gUC9SEkBk2H2K2cQeNG+lvQ4sNKeBOAvX7wltyv69F3JiPF
nEjxU93NOaoXDTGhnsSmmLZzkd3+htO9ksVVuAggzeBhTFYy0xNsaPjfx+L1J73xvkU/3q91QgZM
HiOjTr5rUeXbGIYpOuemZ6Azh+8FXq0Yd82vlGrl8yNFBhQxMDnXSC71QtbF3Iwe1MTDXQ7wkYUW
qPtuQ/nWtVo1mNNQMhBAHvQfZwyk2yWq12QuCP0ee6d13VCPP4oYiaKZgfvwTFEl3hqjssyv1iHc
MCxEmDKqqDNCVquu7neEclRYQb0E/nKYPCdSTBZ3JtqaVKbBowOugkrmke9iBVXp69YKbP9e1uqs
oBhBMMJ+BCIsruBN4O4FTVPOhl3ISGJN9cWW5BGQEwjjxm4SLSQ0zUHQ2iQWuEY667ToHeRBtZBh
4wdtFua6oHuGc5/a7tghSuX7pQbdujef6FnXLyMWFEi7fdejp30Aqk5kcDAQ53RvlrP/rvU+/iKO
wR9B5q2Zc0A5A19XiWCrqmWWD0aqrakaMbVE4kiIRVEq4kpCfROfR6Cp2ebdXEP71DZz8fh2ckbx
QA1UEi96XdFBA/wl7W/BFqPAAJxDOfA0bNOEnWmVhj+2OznD7yYfdUTnLlrxYimqyF/mjReFil3u
14j7G0i4cgfIWk7p2a9SsqODyfVZoa0Nvzrle99bngLlYXfRtY//pJ8UeaXx10vloN0Tleht0y8o
HCJx/MIV1ixvF6nV+xxydzMW/VSnNs7LnoLUVABKqFXnLxQqBzDdU1TkGnQ3N2+G2jVrnTGGUAU1
v3cPJek6lIfob6Um6vywPAmNkiLKCianCdeTLlStkQRN6gCrA1sBV5E0ajdTuMU9Sx7TInPd7jXe
598DI4+F2LLJrpuYEfbgrAXRO/YXLK+nDRlimKVKVYPQ1ahvlGoH7o5DQRFNWqmabFm1BRDxlqOH
i91JTto6sk9T0leDzDnJBSTfgONDIJrLKz24ql3BdW1Ayw3vYGZlLvf0xjo4pS15VhJSnK94G7g0
8ojMP/XtXJHHP0wZZE3/15Rgjmk4GS7w4jiRNFnW5VC/td06ut3dvNM4lGE6WxNkovc1x+2rBWsD
955PdY4n0q4QqjN5JFkER5WClIkv1RAeGjUaU44kpQ9jlXlnh2x/vPwNqPC/iVWKRwuKkEiwS9wN
+HdevzzX4wQliruT8PNNAjkButvkQCUNqTjGeM9wdSKhcOeit8Gd1uY4vbovdL25X88odprRXDVO
KrsiazzYQEue/krV/sAk943Zr51+07Quhd8DMZHxYazdicIQi6eYmAHVdpHFSP/uxU6k2obGYCOR
GXMXxZnfBA8UtwBCtl0LlMlC4+o6qZxwsRP2AnpTe7Uh7GjV/cP+2R/dlo/lw5Ei1CSuNb2jyJEK
0Dmj9fCSSA5g0vp9pEsATTk8f+fIYZMXYA90LKiYs5ti46ngp8dqkGdh+Yi7OCby3hlYs10dj6Pw
QOFl9uFHnZg1Rw1xaBTZBKUlUtYtI+rnZalrq8tzW00Z9VYqX31vmx/0JSSDzswYn1dwfli/+svG
TfRYevXePDCel++9FmDnugz0UB2EC86R+juDCYkPxL2PKWjFQL9xIfoqJ3wtTE4Vquk4QcDTQeNO
JblbDgGxp+UO04FWwB+VsNqdyYmYooOttgzFLtjn4W8YBjcOYiyvmSLzRdAHfday84dwuJ6Cw7yJ
ncr7wUCeanVN/Ej8hW20HJQRyVP1l5jKnUUqAXO8urvoBncKxU5BsBFPhseGYErXm3bSkF2pdpZY
ECKeptlyIq3Wblpbr4FLObflwkFbIQ+DxOenWz8xhR9Hyx2cIci9pmzQAHkuZpz7GlEDnQrPj8b7
wCS0tjnUwws9bzSYjRBl8BnXoSnnFgBGVrNkeNOQNFaIpbN7GElSRfXDFbupExntbt0rXSnApD0N
npczM6/hWqyreEHRW3hwr6XFiOVdyEIfGS9tm4z2IOIdhzYFq1HYm+ST0lon3Lc6Z8hHcRoP2PPc
h3ooTp5E7CSxqkABLNvWGC6P0w14aPD/9YEbwjnpoHRf3YktsF9lIzIPuQaH77/xrGhOFRWLd2XY
aEV56uhqnMtsWiH+op6bKzRvwTYPRSW41U44x/bcRgber6c/1OKmsG4BSbWm7bbWhsZsLyo+whUD
p4peAtSm8pNqGK+hQq8TJjQNVi2pWV0S3F2VCxFpUMPiOd6zYSAntv1xG0SgzqIJDAl6k7itz6uv
Lg+bhid2DTN5agL2QD5Q4VPNzykSWlLaZuFQF1h6rw5rwsGwfEUj/NVTxG/B/gp+PKaAkja8DjkI
MM3RkifWzc6/P/IAldssecz8cqUBuZj057aQl5wQxdas3XI81Anjtij9jU93rQgbh6WZKR9gBJLg
Ug6+Vq9Tbce6NeXNdkLHQeiI/yYw8lC0adMYXFf89iQ3oJUYKInY/8avOR1ckVi0LRdBCY4OCKxX
eoSUQGj+GyVvrf+KGWmiy3681HATF1bb4AVmX8KwM84AIJV/yLA2wH9i1l9NSNYd9uRKJ9w6zhob
l9mZmeTpBRosARoR+gQ3uF2S6gA2BFoUGoQlQrd16q4ZRWPp/7d7m3xkDIkp3yaXj3+jirxy5neD
J21vUpbeiSsNcxVfGn42uKHr1qYu1dfp9NW+RV9SnlWQmKTtLi2wD9MHV12j9oyWxxm81gEH5kE6
ZO6YzYUHveIhuy5tUuboVLcTK9lBOoiPn5aMMsUWPbzj0vvR8Uako2Pdc00bhKAeZnvCTXGdLS99
DotWBuQRH48RKUL9hjEMuLCRagtmSTLl7rYqXa+EPV4Mx9iGAzP4Hct3ZtxmN0yDF1JEz+3nzdhW
iFBJHjNuUk/SFhMlD7EzUfANjycB1/57Sgq2iS2Pn4emE19hMlCTnR3iQ525EnUvddHOZaWcO8o9
/idGuShTgujXm7CMpMudoCLby59WwNtIIGLz/jrjS39HkgDkxTjOtAPtau+pzBeB3ccW4LAWZM6S
kwOL96BF3i1ttO7zvVMwdOsQ5+qksY8pbwrVgFSuDYO0VXZkWHd3slZ/kXXfbvu3HjVQVhgx68ik
FAM3H3857ax0HgMJhsLd2JcE4Bgr411dnZyU76gjTgOU/wuXPCFNFW/whsnyGf+/zBL+ZnYzaP/h
lzmpsEOXK6vNkE2ASPygdLJYmFPUoJV5PNiNl/0TSrGYBsyNprjK/n7SuB439AXCijDGAU4+jeA3
8VV3FsErYeAQBLXxQ15QfvQDsKUoY1LX3vk6Iffg5cvKl/XotbIy+uJCJyddYg5rPC9gjNAciDz6
iAkyDi+RP/CJtpp82seWbVVJQmWJL/EWB5dFU7uonJtpj6v46vLdz3/hul7tjfcK7eKhAaBDQuPa
RG4+xgcTwIRL0GsphQ3jbuKLci2JTrH6CAdCj5fonOijzZdmE3b/w287vCF8hCF8Y9r1rVhb1Qta
k7P/kSPG9r/a4+A0hDhtApAMC9CAWSGMWX06fnt5Fc4vp18Or+61R84JQJG8zCPKmuH1LUCEa6nG
BdqsgDkXGrJuf/azBtBCo/euHIlk+jLSMS0Y/ae6zAnnFXnVaShlfVYIn+WkYJ0bJWOBb4u/OsbE
/mjnh9gZMu9opsHG7u9EIBvI28Uiqxtb7Z2DRmgI/cmsjrCDRFfKDmV3tXtPy9K3HGQkk1K4lYTX
S5loJZdtCcRXLalQ3uxB685wbIBX91AYhF54TJfBzI7UXg9oNnc+E87bMNxtI0Wh+TMlHjhv1grn
grnKqAwVCA3DoArgzJLDN12iGwmocGo0wvahXhogv46j5Hj4Cu8amUGRWH5gAXx5oEhzjZNz35UW
AZd004fW4Dkf6o7EfRQtfxXddwfRwviFo2PIKDptqqEK4/tlskCtUe117pfkA4aGlwso19CnVPCe
dW7IX0PMDw72PSM1DhFdmLd7YDsiNlepOciMKmOY6V//UolYWupUxYlH3Eeb9uDRgm8QqD4kMgHj
hNOZ2uB86oMzdxS1/AbnyuYUSwssxAiF7GTzZdnxAxImykPR4SUw16RVuJNsdi4Cd9hR8RA7NpYL
gNjfI9++DBmUfbb5qIP9SQbRk8o3UUCdNwaLVTkWaQdKGfpqHLGweVBdDsVhJucsPV3fEXxbmLbe
BMsN8zfmy43JMFflDSEeF51kH4Rn4B8EKPl7t6F+MRZG8XoA3rjz8AnPqxou6/YuKidQ9aej2WzT
d8XlRcY0JuiJkBMyukM61n3HykHGf5qoZsjg0bHFYFyZUXdMO7/Op3dpgtHutiAzk1jwb4FXkvLl
SFUUMXwIyBsaqrd5a0JNOQYhzKBemtBA9xWH0MCBVaZ1JtaEEHcqvRLTKs15D3AxkuTmyipomr1D
xM0ra6XfIGvBft16Suajq2jOruEx/5cvd5IRy9lq0rxnkruX2NZ15/JaGFrgug/D4HEKHk5n3Mee
hfPczIxFWtpl33/W85xTW1jck5c5AZmGj7vuvZ7ofAUfzS8jWq70B7MbsfLM79eTeXncPXl1M9r3
KxVPh+fjWZYDYiKMKZBIgD+FqlvLpdoZJ75WdC4TO4lbmM5QFbFeoQgg2X+Cw/rtBU7ztUFvpYVK
C3n97JluhAyY7SOY4A8DR15pCpMcrum5KmSZNW6osytjddoG0n+GE+gUrwltmKz/wHnQWkbVsP9t
7P1wc2AUpqDb35zxFxEKAlWZITu+rSSjNKnyyHwgLyE/UDM7/7bD472zDNs3cBrW/cI94pXxXMQU
ZQSnDVYyMGdzYpr+HnoSNrj4YjgtwBZFq6ZUhv+wxBxal22kjNMy8BRADDBbb+LdwYh/+euFyr+1
Lt/TECPAz7jK+/qhpRDp3K7wmlHJENCR9ZOG36YIS3qRRbOgkesZF59zN4G0pksJGPEIp92S4XLQ
OH+xdcxiwCyzm8RoeuDrjhZaSUx4YIxCeEmHaqMGQcAgQcPwOGyqX4yocwDZ2d7sHYDnvecD7OM9
20mkigoI0fcDL/Xb8cKsp8zG0iEsjKK3NArouohssLvfUT1xfSJbTKCdSRno27b4fV9l2P/RI6lR
+wMqKoe3phrCo4Fyl45XnJZMJeLMgwP8hfxfyMa6MDn4gdyxdWBOgu9MrdwBu76Fi5ZoPFF23GRA
yT8p3bp6AIpkypLX/aGZ2i1JQPeb1duSpBaPXcvRATZAFI/agMk+91GML1yCOcDYKJIFi47aN9gJ
lwRfei4CYaLVe8tx8WcEQgmD/WA+BmjAoe9FmgSYcMx2KdRpPaO07tpuVrG1yX3pLu1v1vTsS0AR
FbmpYd2xrprgWqt/FG5YQVelxSPTk6fWKRKqxe73jJ0IAnMlgcfU0ggcj34dXRjXTdn4sKc18vqZ
P+l3z4J4k96vK22lH8OixfT5qttfEbwr9WTiGxW/+WRXiASZv7yVVooxhiwoIXgZRf6Trr0ydEnh
QGt/Z5JS38zybFK+XVDEniEmbAwA9H9vo/rYVyw0cBNCp/OsqaUKshlQTL50hs9mrn6oZEwhgKJ1
iDTWWQSs2gEdqSZEd+myR8hECMxNZobJgxQ0TtcOLU2kyt4UzI8tFHaUOo4GSMgJFTuT3xsqV6vj
p/XaS5lmKorpWLfS4+FdOqk7ldGW21QGixXUxpWASX74vKiimbtBJ88CAmjtuQMkCMs7+Rf0FQjC
Qeq62PNfuxqtszkh5yu0pfqnrCFylv7cnaHRvg0jSvNfb4X3aFLgBSVHW/hyXXtu1SWWFg1jqMtT
zjhhaHuBpa6t3BFieBa+ykoGh8bIBowrFnFcrJhb2AHnIdxaVCKNygw7AwRW1cF3fsOiRIzReSlr
i3G32GO58WLfVIhv5GxqAt67sA5AIdTTlDm6lzEafM3LLSSn+PV79iGLtHqvFpT2YGGPTIt8RW9w
yIRqQT29BDjeiZvBjxkUCvuGpVUkcy6W3rzAAGm17VahJscWnV9izlP8urQB34MwrtO48/hRBy4u
MtLvekd5hD2SkfR5FOR643Ax7cY8h5iEmAp88rGzRFzsPKs0p1o9EouGGv+dp/GTmVXZVSHMDqT8
youowNyTadg3Cw2AYC6GxuMdXrB3eJnR41Z2nnpRjSwN80bQ4y0DjlqpgvQnfRr+oy5yNH6EOs9Y
XdxMR/ZajoMIdR7ve5ysgo8jK2UkRA8VOkLUfIwjhrzSmnb0L8xxkk26234vM6CyUXRqT2NvXG5M
Kuz9Z4yNcRy7bLGP34hIe+0SdASQLtzNyYuHRp3NsR6t4lDF/VROwVkCTjzf9SWiEQMBdPNxBNo+
hRLP/An7C/9ZFIBYhQodruIk7+hoQw39s8bX4kEkI7EoAHQFuKWh0qWzGvX9LmJGoH+3jsnMO63b
rXURwvI/9dEKoRio9lmLpwxI7tsjfwhIDkTXxckrtKG9gHXSvgHaRuZvTJCF8UPKBvGZc/d01x6h
vqn8CFLT48esKtOGWZFYQEKFjWy39m5lVanHfEvwQXF4wg2eUy7OgPJkWO5tjpH/UZvxI4IT8+bf
KOPIDvMu9s/e4QR2CgBwRk8LwmWng+PqKF0pPtCuP4R45cUq4sMhBZuwNS8SwwFL3yQMLr+kACiV
mTwjxcChhJn8IbVXoJmpx+Zdu/ErTFzRdHt0ETgo3H34xCLIHAZDdGAVgmOhEB0oAbKgRos3acMx
s5Vc3lAjDDobJcgfIZ1yiy0O9VylwzwbFG18wOR1gUgZfhqXaDXiJBN+5hMB+NNvO99RaPAykTsv
el2QRn7csN4wcVHsoRwhaan4bbfC6/rHPLUxmOeMZik5m7KGQQXbtlPZJYSxbCiE+ef2ep3/dPiM
dlcy2nQmkV/9V8IiJYdRKZ6XqTaLXsxpCEnewz/aenJGi5pQ2hAavNyjbvdA95OH3qEsQEwPoDIi
tATPpt+6UbNl+yam5jeJNmLzsZ0okD4tIqqh6RJjkeytMNtNKQVuqQLlf2hVJHT+yvE9BLXNRc6z
NJqJSP+COLTM8tk1vOHVsOWD9U5hzGxQIbWN3LkI8sGSS/8zOEB5McSFzs3QeqyJy+7DMK8BetWo
dcqC0bvZl3Kq0tjP6tPCFWZz519mkIYb0HPqJp8j/O2gBUz0yBQ4ReNcD4CkBxlPhL8vC5VJLXoa
wDdmbWi3g6m2b+/2dDXzT/3Gly7g9o34h6UHefCi2VYrRS191kIFZa7HYsRJr35fH0/j+S4jUbi6
eQnIBMtdRQEo/B9vlaLTOOT+T8Od7ek+bOuvInyGWc6T65GDCQziOQV5BTHeOGsGDUmzklKikIxJ
mJ99KaQs8IL8BsethD1ZNMoqOmaC5S4QzvDM6FP24tQDTxpAQ+EEoJSyLqT1j3QO1eNGHmXBVdxZ
JtXMrBYU0Of9XYpYLU4IIGkoXPeU1r5rIIo7ET8nrULthyvSBvtkicpI+WUcZ1PzBgnblDyUhoPn
bQzhiZD4vgvWNOLd7l5lnXAlFB7Z0JNucMDrHM2XEyx1h4XH+t17Ij7WlSnaYPoQVzJmlscyFq9j
qIgcQ9UJ9OHXiWNCYmfh5uoIQSRrafQPXQdp9blfXJiBFk1jaX2vLZa27XVcLxdWRorDjujHtIR+
RKjv4xQgyfs+cz/9Es6mA9LBArIC+k58J/SRwg+rrCGhhZZWZbLtRX7DAoyUk2vOoz62gbpTzPEd
BKjUKqB/bigUtuneeO/WKh9SEUPfoepKCFF92TTVYtfQ+WjhW4fKuFmY4Ag5pPLaD25I7BtLAPwi
4WI5jhT9Vy/kFSNbbCNojGBM4A3nU5+mU2KoWkuaCyYTU1wpWrWook/zyajQswpgqIdqw8oiq8/5
aRaV4vzG/y/NT/UXp0rahg4QxdBHvAzkyGn6+1C/gw0DizvoMT9gSdBVWGH8azpf5ufl6Z4MJwgz
90w117GfBLUPDcaJiblRNt6x1ysZSAP/Y7rbV74++C2uyXFTxGswYyudLrLawrO0MJlOJEiEJr4B
3rXJn7Mw4VccnP2oFGFej3hVjKQNRB9b/vtnbZig27Mt2fIYU1yQkURlHV6hPxGVSFl0ng+qGYrc
ZSQOnXqCr20ZiAeVgjWiDJaicgSeIagJbLqi6jBZoGxrvn1jY+YW+tja0C6YfBNBjQwGa0IdmmDo
gKgYxXMkKf91VyQ1IZJIQTgYcP6VTT/JKbxhwirHuJeoTLlCTYuBbiLd9sjp4+VgHeygB9RDnsVw
0MZGoD0bj3av8ygpjfyY06PpmLnGEZuMoPydsfb7ATB4EbXvOPJVHMLw1jcYswCVpk17La71nScf
DDHj7KcIHzfAE5KZhM8xXBvRUEZXmGCuKXll35E2rVXDx/Wy1B1XlspG12mYu0QGY7EdQ9rxRPbj
Sf+xA2mavEkkD0W07M4JYAplmWGg5jJNOF1kd0zqWpG24k9OWVzWUEAxXMwPF++KJCkT+Pi5tQgF
1pUkXfAMSeHfRpx1SyiXWMMcUDiYhY0wleN8NYwF6M/y02SCiVUI9947QfaehnTS7zX4lcimQTZa
goosSZEkoc2K4gKVxcgtqFKN2Y0lgY03umi2/UdTYTeN+YcJdPMlnGbj1eozUkrtSWE4L3J+2kUV
3aOmKjwgIvjj8LaF1rZsDtOxINUvmnqYJYfmoDhOcZ7ubXf6Q2T3E1Za28hbPKlE9FPmpNartJL4
19/S7qZv5JcKDyinu0ZW2ATilWMFDTLBlltiyACWSY5xvtMF+UMLltA+o8s0L5Fim91cH39IfIl+
JW5cBnMDTQ/SQflBGrY9NxGECRn6gyJVrfbUg4PUyD3zhxHRCuMzwrcoqt6GhclB51rWaI+FcayC
vrxHMiXJgZ6o5ALlFFEU72C1vRN2qgYBotmgKwHT72J8sCQTMyOEKNltgU9ltnHWIy6TZD2r7KCk
LflHBkMt6YC8Prg7Z13Hy4C8wvWv6TdG3zwUvUx9pdWOMX4M+1HefN3/YGbk1WHVKxpJuYRZw74N
yhWpZDSHcZizuNn13+fE1EpB4OqPO/WqojaIav/rohbzk5kYy+1ar6Qtrs/hDoFmCVsr8T86eBrx
jDEw6mXeoJZ4EvXPqqEEfm5p559myp4YSO4L8yepwXLIM63yTbs3005m8lTIJ/h38d6HmvqYPDVg
xVEhVRdB8RQge2Om2NXeNPGV7C+kQE+YILXa6FHEpwPvbZc9uHiAjPoapv5c8RRJ4UIOt8gyscIG
U1VPqmzPHxlK2aCnwf5l4/bh+iLIFxqtNkyUOlOMF8myVJXovxgocVIbo55l1oBhRVk4VJqrvs41
OlEaEYHp+nToiyXsTSxlwacELzWFM4KAha4kszW3oAqvzkfxZy89aRyHIy6AGPTBgW1IXP1wV635
m+7mT/uag6irTwL9ph1FDBE/dtypdAuFtBDHPq2YDK2pl38ryYGHCJ1RoHYS1XeLyg+EimfDU4DT
SUx1hQ1Ijk0Co4DT2WrnugjCyQuqISeV7OHEcOjt33Q0vQ4lpGiVtX8CQtxsGt0XjsgWzaceP4H2
JQR7UrffBeDLF9joAx1Y17tJxjqncuDRPWcy9un0OKAPDnw4MEu5h6ur6SATzJXj8sPrjOvKx2Aq
O1pkvBOTt4YuNmDUpTb1tHBSBVpUW+mMS2uQG4uZGXws/X59WQUXOHmSm7tpVWQSey3tX8w4TYWB
E0280zLzbvx7TR8Rt2niEQFAFeNGjGoWmzJjZ0ct1tGZ5LxMIQC/oKXcsvPFZeIvMWhzTF6fdAQx
NU28+3R6iU8prdj/eolPhxMrSpi3C4iYhZeL7G/qMOrjlORvl3f58WPLpF3BIljqyKzuWGS6xyQb
vE6m10+qq95bfk/ecqyIWWi/gWIyt6KZdueiRLGLFQWMFQfSc6bdkd1yABXWSbcE0kZZp68IhILJ
5b849GtXgdO0jqSbpZ677rIIQ8IMbleUriGYrpbiiVVRF/dCPIf9WPqKnl8HmGdW2kmrWAOSYya8
RzFBz2WlfGWaYMaUVb9VojgPSjMh4ED4FUMYXI7jBERilqVNkoVHi/xrxpnG0MwX8XG8zUoSPpxX
6UuswcnQ/n1gwe1CP9m45O10QGQxxRiHo0YeoPYbhgk3fLgagd7bDdXDAbbw+X1hOUw3L2vn0Dc9
ODDiZQsJdjrRS8lrVaBvn4xU5ILrfqxoGtkizyqlwL+2iRG5+0kw6iXfkaHzrS/VbciiU9IRut74
vwEE+BCtiDAkFhXqH2AMpKwfqdfRlOsZWUHUYgm42YqmMVKyYBpqpTYWnBrtNS6IjnahnmeouM3g
TjN1ho7LqWGrEeNCYoZl2GPr0fiGKoW4Prn0RZm088Rmq9jlJN0vZTFLTklpS6U5IHWQucUALLnI
PZ6UZPmT7+D/l4iDSoKZ/Ric4W3LRGfFf2s5TQCJGTWADET10SOXzqM21Ya/akLOO99ZD+LDvyNn
KLOZDD8LI584QynDYpBDRQJYyQTOZgLibmyg7LV2pPdTprWSNieOlay2FDZnIQiMTAFiAOqd7KMD
8JGxXyZKH32zA77wsuQY9OJyly6GRH/8IVruABO7XwoNZ8dH+bJwQlDyyDqYdoT33l9atyf3V+DT
MqF3UkZpYnyUgM6xsyc4MfQlu+eeJolWh/DAIGJczqyRJhEOxlwlgiG9q5/hSsGsF3ika+tN2RJI
cIcOGSKi45goO4Uk3HGet1e8/qHKTu6an72Vk9FVmzOlZh+YC4aeTsOPL3w2v6WSUptMLmZw9AXV
I6o+1mNIqrH2v8ndDuaemDDffDGRNlKs018E0wTM0kl/KdRCPhJ3rmJZ+XoHMEL2qo00HPt/VgFi
2dZ7b90/iV1Km83rP9aLynuGpOZYs/ECf1zN89edIbZTXQ7B1IHHKcUrUzylJbdV9rGYJ9rSftXn
QpK4+IwJNvp/H3dTs69YYh1EUB6mO6IeUKpbVdRYT6xQXkH/aexbrkzSWMPcy/w1JsFWKiWW1N4Q
gqxvxTU+2YwbqWnz1hplQS80+sYt0HomjdlfqrE+P6pC05BDnsYvn/VWsI8v/BTEcnfPkFj3WidK
9Bav4y9SwQXau5jqnTiahhX1jD3B5fhjvP0Bnf2dQt9EzHCsrKRxg79wk95NwMTJVtbHBJAOLzvm
BtEcJ1YiFs0YCVY7P55XXhU7HhHvsXmRsRdgE+PegSpTOG3Vq/jZPBDGSE4YXDMTwmKdYZ32kK5n
JfxIadvzbUEU36P/3K0Zv/xWHV0TP0Lh3rs2yhCZtCsNtKVBpEBEVNFFtGJZsCKawdsDffc4svP4
+wgL6aKFgZqgIfP+s9zQaTsM0uH758dIpCTLshmh2OwOUAXTiS7voi5ccNqn84GXMAh7/WIP4Apy
O1WTZtkuvZbLqi2Y6w/G+aNoXIXRSJCjgtltf7gpOILh+KQZEkzBddntyHJIdVcEtCPUyjtrcEW5
HHgdPCgoEpJIwWfw9B+zToQxr33B4XfluBG6WMYMYxfz0Ojqn8HVnLlUvxvHjkA/FuFcwF23bXIx
O9TP8IqP7rvWxzn9mzhDCBtR6EUDqA4fMMNxMELcSpiwVw0t69A0YLMjxJmpOzQq4wC1+UpMnjYo
ll3ECNlR4xSbyn52EPYzGFrRHFHQ2Jkf+vHDR9S6ZDZpWXu/f+QwbJ8fv69QSlmT7G5btsrxdmk1
0Kz4WBvzqq2604wV5m/XO6us4dDvyMCxQsTBjI1wvm0B2TQ+OyJrXNRqpLSa6dGtLnDIq5vaaVSH
QAsWAfZqV+SqGhmMQIg7Nfb82MhWiXc1W60Fi6QY8lB8nLMjSqb8qPzpZgvN1NnBRgf2Zt5ZnIlI
/SKjEfAbpzk7Hd12Up/FBYm7c531LLDXEVz0jbbTtSooO7P/epuqvoR2EdWTMnjR7EsHE0NMvZ1h
KJO4sMzK+CI0hdRlBytijEjAyQf7afXzMBk7appCUQ7+hwRw6jDNXHmQoqaJmHZ5R5w6lLDvCZ/m
N13Hiub6jqnqs1k5paMrEwHlD7tbpHfQhXH44kvejTHjqlvTiSxCkRn0FH59ZOPL3hyfyE6EfvRi
O1HqbhTXxwg+cRW0DYjjK/tg+8BNj+4r4G3zI1W2qq8VaqjlBejmDObRFO7fx43qKwKiRqqQu/Yw
iYu4rGaZ8O6prH9NiwlRGrGrzkAv3P3fEXb/jIOA36J4tlTrC1zArZAV9AogYg0OP9dFt35bReh6
pqrupvYySS1Tn1kxzGs2eU56oea/TJlObrOM1ESCRtW76kriJPz+gITR6ZK6pL8B43JV5C1wPT+X
9/otDA9q6jzfuc171ReEJPRnPm4/6oi8msPLrpCgN1YRSzgTyUQFslgcnU/n7wpy1+7A7VnM+hdE
LRKWr56paqQ7Qe7+wW8dr/w2+4XVPWSUclQFRdSMwb8IAJhRsqL3Y2nNfKrEU5OA8qePuTUTj8Ni
9ReiAnJzuQZPevyGzkhqZDa6xQkJXMkPLLSJjoDN2+infd1BNbeGKwpG+6ffR33rrUvAUiwigPW8
6wS1KND2TGycfl9J3XvcIMS7WobLH2SIGH/PphjGf7glw/1D9b/nBRkK3cS7jtH9fubAoJxaqbs8
+2XKBuyCUeMo86l6kE0nq9aTWrSwKfTzpcCfxyJi7t9OFRUGUZ4oLxelMrsYKhVIDoX5r1Iuupg5
Xw/lIzwaWsbjoCXeTOJmOF+xOlQRwlQZosExJvf0vS6SSRMwfDsotNjdP4OBGKPpaSw6kEgq8us+
GrCdilmD2mlodTmRtMX+4I5JbShO2oi0yDPIS23rc1h78WO248idGaqEXGEsZYnAx3DnV8NGGsMJ
xO+Ru1pNBy3GoeFVgbIQAOSfBkvbNn2GpMZ5a/+xRy4HQmeml6TgEG6eqaBnTY161fyRHfejE6Je
2Eu3kRu532Nl2O+c0XL2WrOO3+HDurO0+qknD5LlUHGjglC9/N16NqTYIhgwF3DxI+RDgaiOXTya
o/Cdxuv2SE3LNw5wLOZxP6N+HutNDugnF6Gzp/HOpu2vEWdtYgrRg/KpAWWuOCkaBo62TSN+rkus
eB19r5KmvioQC1C67J3KqvtmVDUsgZSg7Y8mlsCzWnJcQizSqJG/iVWAGDeu+2zjnvV/+zpauATD
cwPmqehWVswQqiBBl5t6zwzKJYqPRB9YNUsDSw1vWoVNR+HyQV1ESXupw/D3w0qKM2QVoYyfMYNg
EP8pJeLRur5Imatvi4vPaZrC/ZHCwFSuKmo2TN2UtqEHw8qFDq97kD+BMvWTSoIBIBr77bGiIUPj
vWnrbjRbozUvycK/5d1bGGQd/Rn2U7ADDgzyIwU/ApjMherjx0pOZxkNH7T/eujrFrhkO5yNW0bd
CvzP0CTDXrmyY7ryuuEjMXIlnBnKkXDPAF0F0mlGzhVaj1p9cjLjW+iEAvigVj7B38AdjzdbL/AV
FKV6EvcVb6IPojAcXpwyIJFcYDqWIU83lQ/cdFzWfmYtQ3BsFbNPPJa3PyrA5jlLoBidBy0tU3fj
Y/GPX+vcy089qhV64Ll32ywNm+qwBJLS2M4qzBqSKiZsJ5Gip4MkCf0ydAaMZsYE5wzQHB8qqmAH
lUcmgnREVxBx4dM2vH4rR4oBAUyuY7jF/DhVZWZfiVxjFnqcDvwH0lVLHhm2SzN6Am1YRSmpp5QS
azRu/+fYTzA4WfFE1KgAkDjZR1mwLTpexSxjMuQNv1Z1XpaM5l1R4s4KVjzZ6d4Y+h0wq0mB/apE
ba+my8rNHqDu31WivYNXiknKSezIrPGpPZpylC8FiF5KLtEwshWNnXGJP5PHUId3pN18QN28ZBJU
IPXMxxPBEYoINS+hOIgstPph4aaZvwvNayV4bimAIaN/231ppZOsypfDfwzdjG4HGT9ZxWdRbxgn
qIoul/AB7uJ7BqZDC+n/1rTTpdVIzapowXWzUevAUm42+Aaad7o6a7wmZxbcNDrEDXYwW5xXvJm1
Mo+qcAHRBMg62edgPMm1nHv+Fo3VaMggLA5RKUWjmvuOKQyxUkKa4fPJt+YZLwR+jCjabf3BFbXu
y6oMJWmySEPX8BxG+zJEyiB/oFGy1JWRnP9nLbTJFDpwO+esT15GGsqgod8atOh58GWNS9iB3wf8
ehP2ILlFXEF6Ry7VmhmF2JNn/rWrEzmO4+madJsPSm2XoxjMF/grG908CNlf5ifmw/HM8k/QaT08
yIql44tT4E5XYVgjN8lVRkfOaLqUdz4+aEPLLZKPgr+TLIhqyVQPnqxOYbm26qnkeqnqjAkB07Gt
fZ2cW8AfQVuvpjYA87pA6wsm1GlEnGPy7bj4yeaLSl8Yh+6FyUv/l1jf3AJBkWEDoD6IPjr6gzJ6
1hB/P7tawOtAwW0aX1llADOx6Z+uzWe+6cMkR6iFPfi9jkhparl2ty86tud0dhNBvF8Xgcz/BDOB
rX/D5cLBdOcDU7X7ocnE/JCe1983allWv9zTulnogefk1D46AVAiNJTwWvfwCe+zKqgWjNpQx1c+
tDES57prKAh0e6mcUWLOfjTkz1BApKUujlWKViTz5/a7VSnxklSOX/BvhEp00cX42lOFRPxj8QIr
j6b/1i+4+yHP1yY0AAHJIVsD0umVyT2EKN2pGxQOOH/0X7Zdg4gxiKSeiKjz5QU/ezIfdr1ozynL
JV3ILB4byEKOAreo4lukjzS7b31lomgppsi6JCwQ0qOgSTa3M4A/ePHvE+ge4+5MPM1DgU8tstx/
sWk9IPEPpr7WlbobGKFrCeMpUYgJHO9woAEEkCNPn7KNlJjyNU3JmZTV6esyWaOKENPySfNuDEns
HxE5/PzfbBVJtFY7qzfw0pkm+2LKEQrcwPVj4ts57G4xyDPhiI2xJOcB/2dOWgecGGq1FnjtbuI3
GwLWmu0X+Z8++XTrW9Lkyx0BV5YJ+9E/SN4ActAq8VA52vf9nSDTktG4fnP4HULIzNx1omBF0UUm
08Nh7BCjsh3VhQ3qn52cTdtH4aJ35NOIobZAbI9jRcsXFm5qTvkKr/KdgSX9YDOHDqnc1dQ6iqmj
NU00t7p3gR+6S6ey16w1p3zulZj91O7ny5FQrGTQJVpbSNlKbqX6+lb/s9GD9IKbyMz+7vJoXmlB
mFei5nJaXBVp2XlEDpIe0dBWj2J56TMQ8qVFfv9KVLHQkXA2Mb7yM1ltCQRBz2NPd0dfFMqG2vSM
mCDpYlixKhzpVpIUowiL1HwGttVEXjHp7PJHfDuFdDEt+zl+hWpF7Po7hdFeMBkezNcWRjEtvK4Z
uE4Wki0051st6fnBFrIH9GQf6vmktUc362w43RaNRkXt53VB9DA4zeuqGGio7Srt75mvM6f43S8s
yB8q/LvLyY/sFBF1Oli54m96Bbl2zC8XeBOdqhAR/lHwu+sRJRm6VtJe2v9kxc3tlfRYbJxaKG55
NAkg9kgFCgL8aGgS34Bn6nGBf8ZfmobEcCm3IM3tNJP0CPMaO0mWaaxNE4O/zMpmwP5MBClaSYXi
WOmSt+h6ejE/xQIZhAZSM+oZba9UJkvbSn3f587Gj/IL9cdPkuRo4uXBtdP3h6JorpkvR2nWNGyL
AaHKTx5fIW08wHUbweQzdih1fQftr0pFii7FQ6TtiGCig8fF8o8BfqT3nn2xd9htNGE5pzHPJVQo
srs1pB+pSnnfS+XC1gU1Pkb17SaQg1L4RoXF4NJ7K6Av8+z9G5UZbB/at9A99+sB9/ubGgZvWj0M
9H7CxT2AnH6JbFQcRwVDPoN2EGExvtiv1fIAInWKWOHpODKShMnDDtRRkKyRIo1uPluDkif0ns/l
C3ybSFGZGyZS8v9MAfRR8meFNJf3k+yT8+XM+9C2ByTHcuT8PmWkRIQEyS4RFyC8DgibZAvUsb5i
3Ihl/IGtWbZb+fQn1swJur8h20uBtCO1Umoo66kjRvviP+KXj60Zc6j3NxzGQrwLZTUW/oVtmjhs
EEEt044g5xu2igpEnzt4KdY/+Adg3wiXdTkGRMpH64c7hjWj22fiyg/anJ8NWScCMRHzjFAEDQ6M
0L/aBUCMDaQagK+0SecFctFMT+UG7Rb1Sk6GgAQFpZhhAY3tOAjtx6JZK4+oKG3VvzDWtHogoOhw
Alczx47d/CHvwgwEBEBE9AS30eXaQ6hlPHumF1nwZs5xP0aXsvfMAtAKGGAdCB7i0vCBjnxcXwYN
sDqfdVeXBiJaiNK3CsBtGc38qiGzpJSXURxwgY6F21K+ipQ6WI0gl7iGFP7AGhJ4nFyc2cLRlvEh
KtQz/sp6u6f49Z5s4pBO6h+jMq7iAWWrWZkHRzu7MVRYfCIqKL1oBTfNSBPFPiVDXkI9WFK7kxfY
og6mvfDseBlNRMONY7527zmPMAVTEmtN9gBo7KlSOefFdWxWMtVRFhrCvNTR06ItBSl36Fm/muZh
jqZgvj6/JDfPPikm/6iQiDGodKCoO+yMR0V9Ty6a6tIk03fVmjHAW0auLGT7hVr31qQAUsWr0v2X
TuCdG2ObH+AYNb8Idrie4n5ywduWpJwysUVRmP+9CeojHP+MH9XxDzGMN2ft/0y9yizOtilzCLrB
ekelJgB8gfhDJ+SYMlZ+xcIGcEKV1NCq0Sy2yO/yHsGdupf6QE4uHaZBHiYySzI+Tmf6Q6ucWXQZ
eyHvAXhl7BtB9+/QvMNXICc4OMH8T9fIRqbtr5kgRxl6e9ru6HoMY7MzMSLxxR+YM1ryOTqMo1gN
gXK4aovj5aDATGDs1JWV3BIRkaZRvuGv3bh+XSfWeP5Aql+kki/VUYMix4plos+1lko8aCtKt3UQ
5VAzDXqZwt/tguFDk66uCn3fNfyPxXiwQajm7PEub/iuO5Pjepj8gZ9O4MtJPMKGZcb/dOsKJ5oW
pS1FA8zpTAIxhauXHVjp6Dl8S68g/Dnx1CdXAxdQeNxhh4O3ApXnnJAJ4sp03Qve2M5o1EtyQzb/
34Z0oxaseGsBi0Iei1bPZSuFy4yZTbNr8NDhE9TjelA620MNgFRWBLHQ4vmJqKYL0Hp1abORujFf
Se8LH6u9MUZjXQr31XIsHjoDcz1kqqZC5eP1UsShcVhHmeB1c7k9NhrJR31rNB4Po1Vf5ynreB+s
f4ZtIiosnOTk1F7sE9x08ynOWL3k+LgouIcSxHIsRJcoZ4fO2tr/kdUPBKu8T5eaewCdNLVP2ipr
l4uOgHJ7xV1V0UPsJDIEpILnfD8LhHzgszlA/K55qRKfcyvavxWDbABv6yBu6rzUS2c5giTQAd8m
WRFJZUHiZ3tzq6dKadbkhf3U+qCAjsa8k9EINAmPjvfqTdhsDoBd0OErUAUaUjilzIEiIYzoT7C/
0/aUE5iz6uagTCKQhjquNKZ+jJsD1HthPFu2Fq5Ye1EO9pBkmak1YVJpZGn8n0jdTOFeOKd9HnnX
dzjvdxxnmddb9IuIfvL/eceuvxcyxsRJws/bRPbkWG97fP+EQz5CnHGd2FwyIl0/ZG6G2Qns4dvu
m408KQjwC88NzS8A5I5PTKefPQefLIzlvCgKlEcmt93LfMEQL+3yMKDwg1C872UW6U6Fx0QfgbcS
IYH8vkcstzhXwDejSOx/L3tgIdpQeyXKXWeCFHKFBIl7KOtBvSay//dMKO5RxzWSvfZZ8dkBbbX6
AkaZVIo+xGhtEeIgj70jBSkhvW/otAKK11nWSGJh5PbZGLfOmq3cn2VZNi4/8TopFMLBkBoBbrap
pozNmk23vOLkaUGDnAOtduwygaW7OE6Ds7t2mpeXeNCi6MmvJjvWLDV+2N6QCfPWRjWYj8ft48Re
9te38e1SloclgST9OD9XK6FSd+1OMhvbFXKTwz0quEHqGGDRN+1T0ic5UrPC0wzi1pZ4AxD/2imp
Eg5atLJ8iZuhqFwyqd8rceata3jpPMNNqVenNTHF5qaN23HdjlwSdIrOkbU+5Lqey0ybEkeB6Usx
TgyMp8UhtfGRZZYVQ6LJ6tHDjMNG4gaGcprHgkUWwnnwFKchBo9TiEHHMesM4g3EHCNOJL7Xrcee
W9v++jZLQb7HgRDOpptX1dU2gwBYdsiRgqlq8zpoa9k2Fi9eYN3llMoxvzHYGnOFK8ihVoj7Rhzk
XSgSx0zSIjpV+dhHps2VC/FRFXBPKjArPO9u4ToJ/asiNe+fpuc+w4tnv6h4i9U9hHfzKF019dAU
2b2hHKtTI2rErf/OXKtc8akmP6P5LIEKzl0nSN/54x6su1oY9BNLAjddqBIm7n5Ge1Xj8Lh5uN2A
e0nsu93R2H4zbDpQDU6yMoUfklOb8Lacc82bGjeCKqOX846ye0Y09Pv1RDUxCoZrALvHnWEXv59c
dfqOR1D4GRmVpLWf2uv8mv5kMB0OK5jXg7GLmcbc3USCP/r7+bAe+n7O4T7V0Ny5Fx2h9b+h+ciD
bL4b+BmFVzk0U4mo+QjZozijrktV59vNJJec3/Bb0ehXDFnnByo3i0iUkMQ2zuREZCRESCLo5wSg
nfnQyOMm+jdpXTgQT78jclVOCypkHkpQq7eUv5x4jvMdyQpKWTNBM3vIC0Pe2a0q7USdkXKhz6/q
M9gIAfA0LFD3dsb84Qm2RAe/lMsI2CCZY4sfDiPawVNfhmT4s29bFB3kcfJpxaJN6a7yO2wXhBLj
MmH00Wv97rK8MhtHR1o7YIGqENvtDXI7Bk9Uqthv9Km2ZIE4R4Tw6Z4YbMpc2Rj9YE6ueRe6Woys
99onWI5Wm3ne1U5lGNFYYqPqDGrnUp3PZDJ1BDl8SjFHVqdKPYT+e1cmjs+3dJAOQytynsDdMzCs
GVyglfQlKzDyhHVZIjaDR1dly3EiVfCa11Ql/ulrJzi7PQEAkKuRkcxu2EIpU2Q8kHCZYqE58ieK
EuPEI38z/1MBsi7iiu/9nGacY+gKLVim8QWg9twox3Gty0WAev7582sHRVVILR2TYd0lS6G45EJP
ST3HytQqbeYNUz3BseyVdVu3vHqjEhvM/8XXx0H+pPXHHZ3kgoBNu9MIwbWSz/eUiCa24q9N2Szo
sJj3zNzDZqRDCAhco/lN3xcvugEcnRfmomSWeyQarcukOSVr42a2cp03lc9F/vmPgiXaJTQ6C6hY
zO8VHy96VhUTRUAC+xLMK0rOWD0+NSoZjQPDeURj5z7imGayhAhqpqicdhyeONcjmHqxjJXyzDGo
YrU20ojd0E3JiDRNggPHaSZM/8mnB1+VjvE+jns+55nE5ZEu35+cyXK2sh1VNCUGsbbd2LNlW678
6dKTG8+UCZnq5AhTWJiH02mGqoxDd7j2MQ2NiZXjEQyejgO8nMT6TbOAUZOJ698Q1HW+hBcIKZU/
aNnUBaDJaDETWSsALwCsP0kOix28csg9lrvOFyBDUMwhAlNUkLy0a2suoFmbMRHgZXJ2yPIATcJL
JMvvIVKGeIGKq+8GLTorUeqRE+lO5WseNupS8YZqAFLe/pgKc9IX2176dzWXsJP1/vOM8DFogfe2
m7HVqyR896arI5JkXqfJf8WRBA3FOGFUsGvuRWWq2TwrsuPX8BWAN3Wna+S5FTzY58SquV1uEmLH
L4qaXI/M9hWO/wIiBuR1h/t/rxWsMMCp1O+7pZa2eDy40U7yVGVr5tVSGByF20MZh1qX8OIyJ0k1
4jsp2v4l9mQ30K30gseLS8mLAnZTh++Fk61YbjqaoWpc+B1lL06EHBGxvuffIRUJQukCILvhUse5
FQsTV2t+XLAO2TrxrNrqGUPU/3jPvFScPTndNUMr5UOJwTpUhOckUijdMhgOZx9bkZ1Q4jAs8shP
2Zb0WiSgc/wfyH3L1ntgyQLXcQsLm57RybK4NYYZ2A+Zfy5JJquZET6QkxFHGzwt2ESrOegGJE1G
iO3gajMR9EqfKor/0XY2fi5YrCvxJ/Eo6LQLnNIGRaApFrpR7jVzyGE048Fk2so0g10/DyCm250m
/5nLNVxBd49Jaebw4kQqAV8wdBhy5LqWQzvN0+4g59dUGLuxkrHAC8sM1uyWL/iF3fKTipA7oOIU
IkUCnxcaB8tw1Mcg2d70pbf2c/2xZt3OeW3lFMIk6Qk2qsfY6cHyjCKQeBdYJ4/rDVUMjaa8IkBZ
UGrH3f4WZm4/sOl/OaiwUbnJXDzhfv9nqhueAA7pgphjihysztzrJWpWnw92mBhSN+DNNT27Cx4O
ubmiPm+jsShdIFqAd7hCcHje+v474BSmSVXENeiW10Rt5qfstPHebCQtjBN5cVEWUaOjb/afD545
3iTWHwe1NGLGVi+vtyH3xE/a5jF2ATFQuQiHDlQtiJle26owb3zbeGvXMcKorJC0KCTC0kVWy/2D
W9qzfXQY9a+DUFHlQMJ0pinrzgNme2EMWnV30V4WXVDWyWYnGPr83e2gOGzXxUwyp5obdQ+9Jg7I
iJ7pkZ3xp4SM5ITYfuU6VeB5i1Zuw8aBdSu+8HU2hZfKB0L0knwlN6rbkuCNiAtewHCG2WkSiBKl
imZgm6dvexxVh1/XoI3Esz5oKrD41JeFbYovPcp74Cdzb7CEUc2qOFLdMOpxGtQQR0pjJ/ask8AF
lh6unxHW+SmnGjyret3wCG1lKgP7w/FoHZ/vCg2tYPUg3cQ03Yh+o+rO8dNWA5/2ZdzIED/ufRDq
2AaORI2K9EikUDe6kbytdSfN8ZdzyzFthtDb5FZr1dvQHJGOGamoOVWd/sMnp+bK8B2ULuohUZU1
Smwm6AdV7dPxBypWtOuFBeJwB+YOEltb613lrodqncSCpa6M4y6oUxynOkVtzsNJZ7vyaYz3sHj1
JSSsVKf8woKAW3fQyqClFNSHYGWC6bwVGTxSLBqCSBrpKoPEJfiAW4EdMD7onZR4VQ269dL1ynzq
OTmP6a2i2pkUpZbM6R9RSi45TtDAzWSsl1GWENX/0jdwf7E3Pm62wh/J+ilHA7UxP1tM0D6tD/7F
li8wLZvdcNf4XTHjTqtaZCgdqMR/sk7wQjYSoQISRn1SE/ZkRmILaV5zRNIODaJXJUFqCeIWpnS2
Wnve6Mw6iKFd0scbzcUuyBDFQnmxBlk/apbhe+9w/ek+sVdkz1z5jbpzY9OJ/kCOF5CGkkT3qq2v
otqZEEh/XYvwHusESb/EoHLD/ZQ+7f0bfaQL12LZEiHvmoUORxSW17bzy064A/0cg9QLyO6uMfaY
nsgzAR2BZNvkTus8y8DnH/Qw/h7h1qZpcwOWpHC2bv3aWF9oFDoRfs/67zXLom/rZ4a4Jg9WKE5Q
c9rLjzvKEUauBL2o3lWNVLCfnubsupk0NRNE1xqFCs09sKLYvnEQb1xrzAzw+cTMIfGEjTcJVvTa
MhKHt2EOmBsCVMpVEnCJHnx9cfRrCGZVs4ctizYd3roeomeBI09q/PnpEsGAqMGhtm3uR5IzB7V2
3CDycSh9/7/+yGwplEP3r00QDBWl2yMrp9+ehHwbdRvhmFlwBVv7fXzMZhN+YOqFsAa4CpXzXjqu
mrMl7k3KN/iqYXiGCX7z0pWghzDU8+VowO0hlTikegAVyOJkfFXHQKL5yVLwPX6eT0gbRpmcpIso
Q/9hZI6quWNXBihAmFAcGjIhyoB2qa93050kXxRt1ingwL+l0LmzGl8xP86NtaAMMCubOc85pg0N
gU9RpP5AwZDYz8Qe2TpFxqRlvM5l/gmkNFMM4Zcz8BfxmTOESraxxC+2HA8Ax3K94y6n5SvPhLfC
ZpYO3Je3SK2IfgRdxRUfRYr+5reEhGLyJ+NEWVFjgkVeuC2L5azcL71vOoAJd7vuZHr8t5EkzIGU
DY9tAz7foUCHtwdZJ3loiNWSsqfIuNRExccgoQobtf4sKbY6j5xohs1UZfd+/UX2EO2YieySX1CN
Nn2bh78aEGRjeHtDaH//30jZ/8EEpZbMs0M2lLH6yLsm/Sx9cwMXdtFSRAGXJSJ7cU8HOieU/1E6
+2AdHb/CK9IfBOsB80tHxDt2da/z0JM+Wpv7FAgQcCYxwZdNrfld+DOv5q+sJNLbJhqSofAFHm46
wfLJhQ3Ms0FEPwXbF6C4RMSJegWTDtmM4TPcnzp47h3qwtb/TecE+CY0hd3JfvAlqEzAxyIKw4HW
ertZBwQ25YUGVFG+2n+ebz8Ker5rDaCTL5FYkDgczyGwWw1OCYX5HRmftmll9XhWw+RmprY+NUfy
E1qtPVeaFOO1ygRY/b8rIwKswdI4Ah1BF7ICKD04U2wEzyIqiSoOd0i5hAkk8P2nFwJ9GxzvHg5e
E03pnIjQ5/YTVVStR+C/R1eZKQVoYZcOo3TVsotnw9ViJ72yLoB+pttyxdLN06vVLo+U/BWtIFHc
Lf3uDr8b0pvaclkMRuxpIU9Dm9Ib+sBuqCmgP48SL6r7LCuH6mDIfwqLTLe7IS9hRiNvTtLK27nY
IpTrFksnh3+iYOrliHurPa3stPOwWQqbfFFAn4rnp2ZLXl0Q1s9IkVTKqhx2U5sVaIzCz2AEhCkz
4EbPKNjalY+pXhCNA+K/ey40h/8ukMvY2owhc15m0XSa3aegvwphUC9/aNJMdIfxopxvtLHTfBcY
s0UXvWfoe14hiXj3FEQLLp9p0udRcbVufUHgqODPpgoe34pzGd+zL/V/thayZPGu6t9OAVLhhzL/
De2nalnostvWBBgFmXvhedrcN2H85VPb3FRk9NcWYgUIzs3Kd0Qn0Z2RYrLtpJI/QQwSPwKWxgaP
5g1sKIwkZo/NeMuNDi2lOaWKzU1H6Tbhi/B6Aoqw+yZzHR5zwOPEne4r0Hyvt87nPJV+22u0bkmA
bb/jtrTGYBxeHhrMHBDv7ay97rsY3Kghf9beSEsukC+PBrF6n2oU1Sa3NjZPKyhiMpoClNf6Vxuy
QiY/QH00YHEQeMDd1uWxQEGjrEGUfUR8EZQM9FXSMv4JvXL09ErwnniPH/+eHz6d45H0OWJgvR7c
jl+TIQMQcugu4DaOkdT0yzXMZQIcexhT+z3O+4B1NnTvWU5owgm5B4wQQ/GIXoieu4V/f/D0/e/U
+USUAvqC0q0P1708/l08AFOClXvLG9rKMrOyvAODZd/iaCJQArlB2xP12pip+8NB4cAH06uyLimE
PoJpeerbUPJv0blAK9ppTI6mEJvZ7cwo7DTo+7AVi/e+NZJJnYmwuwX9Mcjs2s8j6Y6GVkkt8sir
9EDrIKbaAKFfHfyR3G/q3Sn7EnwxThCorgCSgUBcZ4uOgCtuOwnqRlcHwgel+3QDB2UFar+xhJ8M
oUXW+tP/IrxxJ5mSnesUpx7gaGjRZ8SXAozermm922NCgsP9qEaBSVuzroSJp+WiY9R8M97sIjaw
JPJ8XhO4OpXsnatfMNdmajrjNw7NxshJxdX8BeN9zqqCWYfX2i90l7aABTdDKyUg7dM0lfPFqLl/
OD47XZLR5rhfecMyGRdCqkF2ZRLVDQc+PS/gXXDBW8YH1uxznHGaZj/RGn1Q1WJdRJen9jcMWJi+
5BMxRV8RIlvXFnSwnMhNGVgpqeliLg8oiQG0vwUMJuvd8a792onnY6GJG4RLZGKsYWm93P5G75xb
RzU6jKAPf96DV0h3PThh0HItJ6ZLR9gES/Wmlih4Dc4XwQZnNPyQb57sHdlNt6ExeVqaYMz4YKlr
HJ1Lok3yEqiNKvbDMaurHnDL4D4ZI638FwAarX4d/2RzGDoslOgX2DbKUJPzHb+GWU8Xyb0oRk40
Rs2Nsitdkra4GBSAKyLHrMTBKx49Jzkd3V+YOt7mhQXoOYXVzlTfzqLjLQ5aVVtbIR6JzU/DQw6Y
FCqHDp1qK1r33prX620Lwu8N2afHrZJE+d+1j7lpJCrJv4NxX00xu73KpNsNR0BFyW4or/nG73Uv
TuAu0ZtOC0ErgD/GwwATkjLgnokrk3IgST0GOUYZkIZK1Fg7g64+KwMXl19YVla2A/neI/0AvpBZ
Vvx66brg7fnQ+g14K3aMrVEr9TZzjGPL5KIKHJc3TECZjs5/WdytgYRfSnhjbrd0skJlFuSCs5fo
rI8fMEPTN6FDi+7jua6HoXqmKuPmMS9HyoNN0gB+SQFWBNg0e92M5Ftt5UwNfCvt34aJOI+81OjI
wIPQsOWZZ0+vCEXdFpZUbRv9S36SEgD3O/CANtW0AhH1sMhbEH/Em8gcnuVfZF3x/bjYZ6++zHlF
HJVLM/HRvyVd/6ZdV2GikoJaRVB7RvVqtwC0PoydtmXWd+hnvEQDsWK6ZmU9mMOZptm6dus1u7vc
C54GYWukGLhQFsEr4MoHaBXwI48OGdn1V5nEwJepA3dVx++XHT9VkMg93cz1/D75KuQzel5XTD5t
pYBsugF3OwUYogjAaL7Tb0kVUdSQ8nsRcSwVJX0meLLBwwhZ+fTYnW7ayuvneayA6WhQlOfl5zzv
aHtb5Fvr3gq19/JX8/ojbbcPxYViGQ2djVNUoWK1fIIt2YROdQNHpIed3vrOgKFtDAgv6x2G5KGL
2UJDdtqEPwRNrRvv0pKrK3pYTlxhJxQvA1YPBve4hZ+9zuwqS97fa9mIE5tvslS0LPgyL1zFxxbr
H7EJVsns+4CHjBEiyLPDg5Bs1a7U1wxwx1SlW8yCqNNTz8jHKVVVntV2SVbDN9tGc5troYqTpp+L
2V2U0Xw5D8PnC6gr5VyvV5aqZ8Wa8zrnyqdGzmJXlcyzTsAgmGx+1PKOHTMiVzA45w3IzeX7fde/
BzrTUtyMoKEDGLq/HBJp0JWHWnNDZxWtqd7dqyxMvk18vtTiGxzgb8JqCOe20ukAVBxlLPoFEef0
yhP/KENmUqp1lIpZv6HkiwUgGgGCUIyXKlgE7vqz7o5uRobUoTY02vBWguDJe0aD9PHDbZ6CCdbN
6qwzIKzxlKDXAQ8gpRdNGEetsQX91cjHFs6L7nOUDxtuE4QHqKSaAmJ8KMCOZ+cTOnbH917D6met
Ou9zMGGgLb9Mq6LAaBMGlZhr+W+a+krvZfdj5sOWWU9xoxrfFysuqSpySORAcJ6mKO1WFzM0ocz/
60MluEXEXS8mIhgUusDZ1YV0gJHSx32U1ZsGZ29s+9cvTAyod6HTId7JvxZs2FCyR2dzIzOvONst
W26gIOJlKfhjgo1l314StvHsUiaQd3en8Y7ofs7TZQLhOzQxgkeffikZYeklRbQd2UpgQnGAdvVv
FKrcswDL4ENiB0Ta0yTUXhUuawurE26TmcqwBxI0KAgacJtG9SgUDh2cb0LmvA2tu31DXhIaVK3H
yBb2Vh09JXu735JsCEDtrst3VY7u/mJmvE4jM7KtZ+oLKup+DABQh+cjScoDvKAnyhrd+qh/Kbzh
kcEEDfLc2fOrUDMstZayQervIFSsXK3A0WVL+SOzQpwgSpD73IbonKU/85r38KnfNc1jHchooq6Z
KYuUCCz1tv0fFmbfyjjh0YEzORY+nALdYhiSCZqVe7tUzKRzyt/vd8tmJ+jBq8oYwznZMTlPJqXz
7VyRi0W5MfL443Xn3t5tuaM7p00zWM7bqrzlJNn7/xMfUh2A0tcMMbyBvDd1EUsIvqK3tCvv4Qoi
xZBSAlQ0NusH0B0ung0WZDZOSFWaZ5qeIaTa/Bps25xwFZrwy3RucTsSYhWtwA19WQ8l95pBinPr
176hC59RLYm+KHZFYiXALuvKRfViqS+ntMYf88IWRHxAsYhDgd0FiDpVGpU+0QM6kT93HDI3FTh7
iAFv1panHBH5epJyPgFSW+grd3B6o0gaqKLEJfWRC8iBrd58QWR/jhF3ydRQHFeg7uFXLAjIL1X7
lk/Q/lU+uMCLQJ7sLFAjmaGedLvXcdEQBZJ9RKjCAOdJYvg4nf708tbgDGVlaGrst8HvPw3x8gwd
kccEmw/2OvUUQ1SNSYI8jp0NArVfLvAn+Meh92p8IKTTWsDWW888pVqKXi421I4hVo/MFfH8dA5n
dlC/LPj+Ew9yxUJ+69O4PgDjCnYUzZDOSKQYcAk6a8CrqWZ3gQMS2Ev+YkwwpuJVfvbGJFOTji4C
FJYsncXbLG30tS+tHSFzTKSz/TXGM1n355izikZAHbfjYBk+II2uxoDaTqn0Q2UwUb2Wivg4uZPX
ddDDe7Dbo0kblAPaactd8QAYK19JF9P3RLwoM6S+cWbReBQmkvuLcHr9qCevz7KoaeXllXjgP4Qi
nomVrTHowf3uUdlKEskwfXinYw1jW61V1jAsJ7BTXJflb6lX6c2WtdMf4gYf/BuDkAbGS9nh67Po
ZNGkA55FRU2KUWqaq2uvRAPdAf3jt5awH/CQ651P/TmdxetjtO9T+ZF+J3/50OwCbdm6YLFU81dG
ii0HIIsRD2++JWbd4be12o/f4feZ9HqyqMfmnuJB8lD3bHipxB1F/kle6X54MXZGqe9SXJaXfatP
rkhfFSC4I6KNGuYwlc2TryY6XGVNT0jQP21udVNWgtPkabzWfwlBVDIYHrJec9CUoDd9j0VvVe2S
w42qCcjUUBH6LuEm/6FkeyfxNG5KcjaGmiG88fHZ0+KE97Hez8RMci1FxGhJAdvmDJY27+PL7mSl
hqJP+BZ5n/3zDGerFyCQwXXpW/MVTnUsu35710kMyd07dXD1qcaZWrbDwFkIuJywdHScXwC7FPFJ
F2EXo3b+KaEoobcjj/h/dvlrpF83nI5xwrk19wjq4WaMyNXzwfaRkAl65wi0JF8dFLQMjG+kEWj5
u4aXijqXoF8mUs9x2lgxPsYizsEHAFCnzK4B0i7pnF9+KcXZqzt0nvDKhm/Ksnqbc3ibnBLxviWZ
MqDehk+3jx0BzwVh3qNK8H057tc6XDY6fGaHbCMFkbCNgjvzwWCVMyli0QXbmqgjThgFX4/3Jd5Z
TzZBEL1zdIsWQIV1vp4SvX0/JO4Z2BWaYq3Fyx43uHqvInt9Ps1B6K7O5niFwoj20pimY1FUxi+e
ZEQ7ymVyZspJPHFb9uCfWoyUbJw8k8XUrKzYG6/owLi+8LKwv8PE88t/huuf+fy5+uavc0FBJWJv
1HemZeZlJsWW6kYVNiKG8qnrTKOm1Ux7x70GyYyE6vB7u7mObOYHPbXzPepC+AmY4KcY4epJ3UeS
dG6Wo6+9HC5iul/20KNjFPsrpXuYtSurp0jth81IKhZRn4cfmvCZT81OTvw3yRpyfSIFuSzczYZV
sCMmlE0DbNq6mXHHmtpKxiSYsaPBnVeMfrNvMYfMjyEf6xehxIav1i5+gweq07DWAgnSdEWMG7+w
jfGBxhEUeZt7/Iva19iYBBkmRuvWEjqEikd8qnJjrBymd/yePJlpeFromxcB8kPtrb269LTGOZ+Z
KaEYPoLjCfT9SDHtQpVQUs7Iad/QckmUStGbBqEFVkjnXWG8njLzIwvbyUDlql9xHFtFs42uzMlk
bSBCGp4ope/Fho/S5GaM1pXLfLxPRUIhDVoALb7/5RPBFFl3e6xaAKklop5pxDS/lT3Ol91/nTL7
NdJOwZdHIlM3mWRxEwBzzsz+1bVsk6BigLlYN+R1aTnOvB+Rg4Tffq93HfZlseXyOTjYmnUnpcJU
Zl/UsIGHv2rPv4xYRd4kdpsegbWfgYNyb5h79TtU+LNzdUaws++Tkx4mPkI8Anw7wIvLcUnFsiX6
6YLH/P5C+dwKjSblW9tnJCjcf6uWEz2dIGDS0FBV5b2KzADcjUr/8kZs8eVgbhITIzwsw+rACpah
IhaLS6PHVq5zcFAi1Muu3n5Z6o3EXDnOMItl0FgAGomPdZQl9qsHa+pLhAhcJg61SGwRkFhyTRmd
GdcYlhiXck7w0Bea9yAa9GgfJjItIr+bfila+KG2fVxZjGDwA6pt43bLEc5dQrinaTR6rQwDOocp
4BdiFOHFGXChG0ItTao4kChzK1SxYzKKrjAyA8KD+VqfSTDBc5KP3riBlvalL28vlpIrq7UrJI54
M9/8GBjQJvBydNnsagYvxGgKznOtqHtNOqW6ViV590c1NwJs2lukPeHUPed0rk4r23d4d7imStwu
G0DviS415nuNvd691ctO+7ZsvHbdX+bd5r5QIjk9vHO9/Q9kszL9On7K8Dbycbx78GPlpe7dMJtF
Su8JX8MLx8QHsjrgNh8QdJRXyLrs5FJQ5kCqprZyYDcOVGut8H1/Mx48Wq8Hec7vgFaDAZH4nCj4
DSj13CMBZUlMpo6299sdvjDUz9M7mQJtud27ReB7NXrq
`pragma protect end_protected
