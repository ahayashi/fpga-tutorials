`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
QCeVQ40jluN5SVGG7PLE4pRXlei6liY2Ma2I+tScRGll6jWhkxFah2QXUMXfd3RR488PrE//e609
VB3xaaUfvw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
iTpfY8luMgCN7pK5xb03lBMnWS9k5lfcOHfcxfi7sjpwTwDJ3Bga9DU96sxs6fIkgv6crM0pIu7v
eX3oF+YIBevnmhiogF52kqx+Eg8RiU8QXvxIOO7ayPVtluyxENQTGczSly8chHzbuKHM9wE2Unwg
1IgL/MxnhZ7Cl59u8uM=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SxvMwhxhf01dzdfD2lxgaapXhtk/ObaOLLmTSac+vHSKUtN5W+GHAYLGrZDd3XCgIRPAHiexL+sm
56l9Z0Vx6imcD/0AUgoJbibAdgP/v/jXqMdivt9D8qm8fY5/vOo074heWbmdih1zEh0grNpZn9Tu
RgolxZsFV7Zrke1c388=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gRaJi3MbjPOo2Vp853rk4Ux6wXZ9LewF2mfUTqshgtqpwjZ4sudaWolbo2dOmi1rw2inKsGED6tq
krOayngpyK4obNacSFHxoMp3gtjWxHAUngCa83zRdkWUkLOkI+Vk5Y9KTT3N1bLoj2gOu0GYDPpg
D9djCJZmDVHqK64PwS6kem9gpqDRHbTDmkuGFBXPHAc94QvugJLfLq9rN8SrcAVi3LEwwo+Pd0bP
J2F+YEDbXM6j6TUX2BjoJf17DbXUR65WSAHqLKvWnv6aDJ/HqIPiZagUR75PMAlua9l+XBnLCO3s
kosijf9S/+Esb8iLQEPmPSDOWOWD03b9CN/0RA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
pOHKjbqkxHkzkHiuylOvhJgpS5P20FRtuRhJwOvg8xyG7V/8Q+Q3CmJK2YdXxoL6tluBykksbPzx
Elqa4JBYvmcR+yiB8BGMIWDAShit4CcJuJD3Dy85ghSc70RWDn15VbsTtv4eTwn7BaHmmH2DVD0n
idWVHMzCkUF7Njc3gB7eCQiKA1LYLlb3DGVt7GcrG2J7ylKADPl3VDYUZHHF+lVlEiHrEL0trxZg
9wFN+ZUlKhO/yVCs9vbFMQO7vOZFQEwltQw0/WJezt0Di9OmZoJIr56zQSpBulG0eMS8ZEw6GzkA
ROyin/hyVzV24S9b979YCbYt3GrSHCss9clqJg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
keQ7WgXoY1YL+dIjhzBkeP3hCfJzxkmjG1GzmMDmoeGbgXpwm3cZk8Hgf/Kyqj1YnhJwaGwMasRj
2OFvARIpfnt4GbGbdD6/P7erTiITUaT0YTM570HKOqZJo2Iwt2IyveWre9mOaOy2O0aDzS2aMHtm
xAUErwBfvaACMatzuEwvGh9Jxh9Ehk0REBsZlmH+oBJw5o9xCVh7xn0zoUUShaZg6lIus/Hvlijz
4rZ8LZJCO2oA0vWnV4QFHI6OBECFBocpjl46na7FUyNvBrGdys85TD8QuIAi509wfztPtoVzP3Wb
Eyro6Wwew+Pfk1J2G8FRAltg4IoBAcIT1k2ZSQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135936)
`pragma protect data_block
V9Ce88h7EFf7d0ClvHy6QsMhl0pwcAVnwoYl4xphrRwiP7aC6B8BxXE4sfHuW9E9hRpLz5FHOM+b
6h98fCoyf6W50bsO6cIKOn0tCclcNf73liJ9IHRQQBl5Y0g2hlHp6GMKwcu3s1E/7gxLIDOxCe3P
Idn7nzaypuAAEuvsoGz3uKl1IVAt5EshWIyAou3aTisRQLk2dE/DlaU9USv/4sldDglKAumNatSQ
UslvuiojH2BRcGyKl1LDgAlGgKKTqH+hSqQKlHH1pEdRwx3LefFLZNFn+gq0UKCU1KscOSC+0VtW
V/BZhdhgLzmpVHOCmUuBmYVgbzAAdTjsgIjO8t0ClkEfnRzsg6Hye4XZO0bOXHNwO6gd8xjPQWrU
O9cv5N2/AXW8vierLI6V2e+9irhzNbwuhUD8V1heDTOblaURAe7F8BVjMdXV2JtmiMRmov3XUNR+
/LokTkhWfJYfjRX0sohKJiEudVDvKAMzv42kZqRUq9X39GwUugJD3j+4XRMAhCRmkRyxc/ESreZu
s74Bvj8ymvWqsLNOJSwRZ8/Dx7zO6jrMA8TPsLoPS/GVW1f35MPHTU9oWvsemqfhUewcJlnn93uP
Cpwv8J3eG73y6VjaZgzHmuhi/7ipRbXsUGr6xc/59vtewm8z4aGSpZavkyO26RMvq1YjajJLzPQ2
ZkidjlvVhugvLGaU/YB4xrW1B8A5EpfgT4pAme1cXsgAqDf1psTani2JdpJiro5UF5THlGc4taXa
+JsLdizd7dfGS0HgTUSqR//X4uQd1iS41+gxMBJbaJ1D9TVGT1QNhXOQ2R/uNEdViX8PkFaPTB55
thKo545B8In6efujcIygy7nMSCILzpNe1mn57uFERTKqpbcgfF7dOqZCtmMoQATZGFxw+bMip6FA
tuAxFFMwC2HBVbS3pHXWx5LzgploHlfkRLx7memWJ3aK0SMrLYRThR/Ad6PruZ3Ou8LIcuyJwPk0
MsKWgmRPIYRFdfN49e4OtqYyX+ilhbNxLEQxkhnx4eYLWjLUhE15Fn/S2JHGujhxYTrPmip8rrov
Bz30D1lWzHbrEPkTm7Zj4F7Iy9HPVKHgiTbCpdm6U5kyQrcstbgLDR8s3FVO3mPYM0CSXUG7y5p2
nS9gS+CkXxkZppFeOw/F7KBF6LoA+oLcrvR+zUBJ/j8VPaZG2hNCygeiIfCFp9y81bFcNLc/8yZj
O6eU7qpjZGNSmNe0qot6LMLhh3X6S0dj092r0MHiZZRuLP2owPXO/DlXmgvBepQld/J0NGm9hhS2
loRunnzbpcMQ8TfvYYsDCWe3hjaZtVwD0K3b+bS0ca190EbW+L70+yxo0IyTszD1B1hZaHhlZU1u
mYlGTj8+yPA45q6U41ShuqHbAKJCNwRshF1rPETmi4bNuQV7HomoJHRTKpsjDGnwS3mSaOrPpI/y
ppjoFWA+NNtvWBfyvAgFAOOKcrM5j1zIBXE8OUVqIRyuNLB/2YduNErEGQuiqiWos0YJGce8MY3P
k8RrQRrbXC3Vtaw1OhvnSLMED/6km47Ns5DrVDNIeNLU4HcKODmXb8Pbn2x8xHdrn0Pt8yIzMUo2
FEtr93Tee2prRylkPKur1RyQir5K1NtnqbsNWKJHyxPNRPtlrkjGhNbgaPr39NGTQqnOfW65tBo8
b8eQmLDgj/jnKGdzlE5eengRKdTbi0VILl3Wiy1HLpz2NU5jJZY86SpM22aJygOJolo7w9qcWxYn
fZHNQuvrMH5GztluXaTtk39hxoZnzjBJh1TPaa3XJjMYQfgXwclKn5LgeqXgbIW0X7rWUt5QeBwp
yu9dILZ4/PmyMtSLAfBZmI+pUwu6sDCZ5hIJqlaBhMcm85tlD5Ydsh4QtfgVZtStrMhNE4JicYhb
BvuAdOsR/I86ALXKFjhQb11T4SAgr6uism730PpaE8805Kowe5c7SCGgGK2UVvuSfonZHTUvwsdm
fcvlKF8IOHK6GVEBty5YZmfvJQwYkHRjNQ64/ExOGzev2ER1o/eYMyQgs1AvoXwhOSy6r8gHghJk
ZjNlUBbsHpQGbhcI97k5FGY/IeODztPYlDaphY3nbATe3jdX09P3SbwJv3EFf7Q9ScA8Fd+rKZc0
4hbvd/rKrC7WbpPEvX80whZ/vJZ0uT+Mh3i4mH81rfiD/RzXavaL1Npz5Z4OnOCYhRDMcym5G+fE
8OePor4NNPQKbPl/OFGFstwEPieD7HNn7qIwV2ntVf40c3QHuF4Psx+5bIkQlPwEk7bwkW0yndLz
Hy1T6erNdABpKGNS9KFBbs9BrnYoUWcuhLPoiv3JKAdqVnCu6WmJn2zsx1zOTbExbRBQJjREZQBR
wTpfyxQLS6T7cvK3t01xiszAAtsEPETHofTT3g+tFnX2Dd5umjkWKNJ5ySP3SY3is3pfwO/TW35U
8BBW5KWJ4UoX/d5s0ww97cSlDpB/1cM5Eem5Ctw18Mjc8evZjeVz+wMQNACY/gB4G5rqTIjLNxp8
vrLtbKrnlDpSnbxdv8G+kDebotPArwgmi4czEnMHsshq9ShtNTv55pNRiOkN0VvIqxMn0tOf1Eth
ZQ6jLZAshcrrPcpbubmkWInQOWpbRItBoS7CQhpCfr9thHFLNR46W0a6vAunGe4UuyhnRDK9ZLAG
ccjeNyrpwJYViulovluYBWOhgvVK2Gqd5vbvEHKWfy91wtOGwkEP2CSTTjrHI8krCViYsBRJaI7k
Yh5Zkn4FwsHkW41s+OZZJwEWjwpCmEAsZb2BrXnBFHHQnkhJvknYJX19tRvvm3Ob8UyV+gzVyuRN
z8tLTV3plB56+hJ95qXlNFst2qgJ9XNp14VjWbjKuuIP8jevVEeUctUe5UtOQIZnwkVcgYP6Y1gb
BrvJSCiTYxV/dPdUgThQcrt/RNIoIVMl3FYblmAwTn2uz5dVtMfzTpWZTdvbOnKQwzxzFFgujVHx
2GT8rR/pTQQLD+O2tsz+xpYFVdNpCh7wwCscbypoeQTVLgpJx8Gt0R5CsEAm3gyw9CT+fMRuoaj0
buyx7QQ4NjWKkkYZe2IJNtythD9C/b1xMxZbVY4UffPLyTSloSSG93mzoeoGVhO9NRQj/RWh8pu+
6W9n2PFawXEuLTswCPP06KwwjbVm7xO5EnG/ULoIGt+hf/TwH6HgnGkikikhk2ZZBXTp6lu/n9cW
cuKjq5/XwzuL5Yt/529XaHnydaN1wBsEGHH9AGA045HGQTP0TspoMhOmkVPaO/xPLXR4a0m+/IcQ
dtQbHchncsM6HgQE+ZxdYv9pXxPl/aLLfniGWQ/7rKnTA2naDQagic/d7HREcV9Hj0RWKMxVYxVJ
gvNes++u0DPaP4xUJJwhzgt2Kp44M4tUILPUgne/Id9eNUffwKoIUS1TBm/vKEHh8vCykeRg4gih
0lAQH77uRaxNTnu1eqgM4hLjVMjPhqypwEx2G7wYW5YGpqBEA4YmwhFhNmCWmCWaZXkrYZa9zeE2
xNmb26YDb+npySjPikJMMslJuD0KZeKtfK+CID1HaVyfjaRZvq/O+dlRjgbfleP8KthamvQxIkSV
63P0ugAed03+MoW+JkSloj9xUxEPm9Q3+vqUgX2iohhApxSwC+TYts7GRr4+Vcpy5BeRkWBvXcRJ
eIQLcTZuZ/J8ZWrQ1cBz7pVqw4aNM5PEx1ZOkNUfofQC+0G6B8k8rzO4xeXa3m2SlBmud545Rddq
5p91nCggngTbpQqQUmclZ51dZRO5tm5Gf1dDh9J7OdlpP0yn/2SGS5d7nmhq/gyNFU0bK2+6L8Hm
nt5LV+BkXDtNz3Pqv72mTOvvBLVFdOu1TvWXoRxp8kZaRdyUvw6ZxGUbopoYNRPVsjtTEJnjANUM
Fljt5s6GtxbyqS4RffvoYehGPjgyKzvthG/BWfl7Ku4o/I1kOPt8stfOBYy3/uCtQIK83BFo9yfk
1FwXZ2rVaYFnXi+0Vrb2FHmAFI8CzVhM3LqgG+EjsjYFoBKDt9thG1QZ2hKidNo3X0DH86o71t+P
yD0IjtvwQlST3e/ZUnNXY7vJdoL4RSHr4kQfq+OYQ4Z43/dNC46Urwywji91SrSpo+kL2Ear/jr/
4d39peeslVREB6HLdOEr3nzz45TcB6MpGSSUElr0Rjhg3GA4/xBH8t1Q+PluytM5XxagJGlloELx
KyMt/5zIr0u2O+uvcx02FN7W7Xw4VxgieCz+0FoP6flPx+JYhp84muJEPbaxmT/jiCDPINETOOLn
aI+UNgfwoHPN/MFUGtxV12vg7pT/Du0AuXhaC5Cn9NMuS/JdHA20KuMKgm0nRzqytHxJdqehm6Ib
PHLlAgSOAK5i08Ah5l0fHt1SY1XXtVO09DvE77TS6gRDvey8cyNdb40XI4yXiod4q7wkL0VuCMZy
tPu18wB7NcO1G0jssXPtILjrBzMoFD6W6TAUYpdy5ugQ8xIDMrnczNJ6DSpMKWdE7FghuwxXbAnU
XqH0wyc4H+b/OpyBzPJ4I++Sxo5ckNbcFLHnEVj992EEc/Ye0RYeQLiviX7Q+sjRfka6McUsof3D
T2rw/X8pby3QEfwfUgFCkAGIfa77lwlNjqIc8hR7ttVPIMCv/GvuR3XyajnuhiEb1a4r5Mbj0d8V
CafiPijVDO21Jtqw1DldXWat6iH3Sr55VdHcoyZ33LNKRu01C0NDbOGp4HXNOk2mI80s+VP8qKvE
LLfDh23Wfg6IrwKhyqZ4/cyO7tDiT/BA4jxVncuONreOIE4k2G30EoeiUdqQpGwhkWwqFs9Upe9a
nll7q2P3YJEE0jgVeUPztcU0jhk5Wt033KRSxKdTCyPgKTRj8MtwU+9jB/1Eoa3y4v/hGidBGZx7
XsyDpEQvb8IM+z0b6csLasjF+4BgIlxi6VX1utOOS2dTB3BzgT57D2gm5GKLoFCq+pKP4nROAota
lo8RRRs53zwnxk73YhiayERbNfniXbibmEP5PC/HTEu4oYfUC2P1uP2mSl8CS1O3sH4chc7wNbEm
3t4SccOuIVua8jfhXZEfcLKNoRYhKplrQnvu7o7Gj5D2Z8Mvw2VgAoc5viC4d6TT433I7OfO9gzp
MLXZQ13r7kmnl2ILJYLb1HLa3QO3WQVUeTunBFOOilwnRovm/KTBfLTHlgiPXTelP/y8OUE2xh2H
I9TbwLZ4ueFBldMdvJQKnoMRjmvMHj9DXSz3Wv0jvGroJ9fnqd6+S1Oc6xRJat34kTV+uX2cRMxh
P2kH19FCbzIaMqyFVUWbBN++emlWwYPmgJm+cugMCticyeDEIEe0nlWzVkKzW4IH9OlmP3kBHtte
JJ5KZ+X46a6ukeBnY5KsXiSBUwYGm5fz+pQ4KoK06Zo0VBjhYdyLvBtC3Eth2Q9cn+qksD+xY3y+
faYugjtZW1lcVJaXKSOBwhazPct1jvn/EmmxKDTuM0/1TGwHYWP5TEDQxzho6J66TXPRQsRBqfC+
iX9lDIGx6d6Q7Vbetj260w8dQDjwpmhHCXKVzpqP1ZhktVjEhRRsidVv3gXcGMKnRoHF/NdLJTKj
AZFa72SJ4PhvWRO2peBVev7TwNiZkkV0q+RDxfi0N604tPOgOJAsXiddNQ7mlC17/Mx/yaSuWgRS
3OJx1eJKXRW3YFjsuqzpbU2dfStawZ5jyPlzYTOw1/7XG6PxBWBuD2l3ZBPPn537Ioq00XD3CrjF
JLNQR4ReWedsKPMVWO+NG33/3AKX+xZbnLzBZC2c7P0iStIpzCjA71HTuGTUsFvdjGextG8SHsoh
BWfhJfTLgMsM9+aD/fIAf92xrvGDZ4Dehzw+++dgU8Eb9QvJoH8kLP4awy8qOtDBD8V6mVKz3A8U
0PVgMe/RN9vwVCZCXMZT6hxVw1ULSg5TX3LJg511gDf/Ued1JbzWRe0ak77lKjlpD6iFlKRvPTim
JwucOUtXS2H+8toEs/B6jAmVID4QtV3JpDww5QiEx1zdIiYEqDIFFD0FSfnxQnQLDGjwslrtLW0l
xSSrWADYO50fFP72ZwJMykowCAZPtzhszTGwxO1GpycMz0oa5bizcKMNIbGTJ/r/TqIs8DLTmCxE
Mt+v2vQfZw4X4akHbws13TF5oSQBpuMfcQ7MFz88eycglLcdcoIKov0hBgdGQoODah4vaLS2DA4R
p9hrxoODFH6ANw6tY7JtyPFKdbfOZ8VxpCAaRLinqYHoWFj2ur18ONjVyJ998nVUHxGWp4SoqdMt
TLC6z5hhjbTY7rPpuHFBTq55Mbc/V7JHuRkTjZx7GpJSJC//L7EnIBIP7woAMRCkkaETH7Mclhc+
FPRh7arAP2jLKobys/NCDxGOWnppw3hWFWz1BHxP75XGxZUan3VgUUruT7bOwBcqqlrxxh7NrAus
EpuwXmtCfJZ78GWb8bmUrd9bzIxnSEYzX6M9yfYktMVPPT6KckK4KdlqM72EWJrgy9FX2I+oOeuw
v3ccKy8HQRmvkX/zUfVBu5ErK2h624Eo0pAVvoWl7VVOl9VWfaUXcS1OX6ARUKjqgBN2DmRuFSw3
kCUkC5jq6i5HJG9TdmQ5Hnc26kRAvnxWA6Jve7bbnJ5n4mU5ba9WET+RIuC2cDpDx0W1TOYxHK+5
8HPa5V9r+5lrzWI0N92yh+csX5F1irJsAd24F1putT5ipj4VgPlfQVzz0Jd0Ga8QrhYxz+1KkGLo
1zMv0c+YUxYw76lbMyxHaCYakAYUCEkrwcc/5D6OYEcer5m9G4SKcDtXq0EeU/OwwnEHWWHh08B/
Pi7KkbR2JLLrayzJjPvsE38pHcDwtz0OK4dRR1PBrYUKZX18F9D148XYXpcVp5WInju753zv+raU
onHkAW+9MRP5uWdwl9J8Sy3ZjhVsjMYx+V2y3Gn+wV1CU275Zq5p8xOMMUD4U2C3NvvHL1qteSy/
75uSYrQe1y9i5D2UOvmYHztXS6cfvTr9Ao6ZcEt6LHN3vka+54NTK9aasVe1sBxLCas9aHg0+bcy
3oX2Td58yHQLhTra0YQF5k3C9Yhlum7F7hh3aTXLR4RpEeM8RQc99dn96DA8IxqsINn9mKAydqGI
2iCRV0ff/B4jATdXicivb0GJmWtogvd3aF2Gor+1wpwZ2BNDJ2OjIJB/Yl4sGNhM23BJGG+cm2cF
IsnD4JjdIpFuK5nFf/DVY7E3n+/F6EOkyw//qylm/ofKr5fwPJswt4jLITVyHHEZmDv3ennL7pSm
UpDUb7falAz4Cjno5Gimq6Ra9s0jnzOHXo03Qh0zFhVWPVZq7VoAw7JdqJu7WSq8qKVx8u2AuHak
80CTQmc6uzBNAwBj/FX7jZuAlRbBKwK/SmCIv3vsALP6QJKlUHxIrdVvWdxJojpbsy+AghCNtv0B
+wwfnfiG3IlZCmYrWfhYNQItvl3Idflx4LX/HW+i8gxHGlMuQDUaSpLNgJsSf56kOlOZeyGFvt9K
dDffZohQ9e+zKow4bfI3QNdPDqRYTc8zOM+FnKNS/aSvOAXeskjCgVh8gDtGCW3jBXjdxf2cOQrY
ig22d1UIX3MStpqUNCueqjyRdJkk0mylDdU+S41+iERRYtUHKdBeyhn22vFJNXmNfknZvKXtG0VV
28hPHF6y81c+h0lRx1lQq230kb8ld4fM9wbIlFPQiDMObTiWvkRLUwCzKEsq8tm7YMLJMM3IC+kv
Bepf7l2Da2Z61Jc3k0MO2pTQdrFqEbZ0AHJbMEvfv9GgAtw7HYftdg/dtRSv0tg0gPv2IlyvyiJb
7wqu8KWS2h//J02XK+aFcJmhdx2oXqYE3jqGg/i2Q63cMKgP6GDaqoexTz0d/xXY6J+Xu6GJooJW
YiXwzD2xdzkitEIvNVKJQH2zL+CboaThdxTyezq24nE4k+83PtxxUMF42JANQ7KFuUs3wwhA2GSN
y7Ntf2yxD9c+hRlmSfZ4W5lTljQIEg5tsNkYq31u9v1eoIW6niIcvYOUIqhyKkEBMbGE9eWNRcPp
wUaHUlavkmvq/8XH9/GPUFDEj2MGWKgwo1lq2ED+kTd4OTert+v5AF2mLn6jR2L3MVO9YVS5FqYn
HWuCxTSDno4hIwgp/sI2JpZyCGqOk/cCy6wjaOHPbE3W9dNjLZOBxD92QBLUpp8cOPaxXimbBzdd
OhMT8t47P4Zjo0qUmoQcCXf6kUltHPwvX/Fvt+o+Kv+b23cL+XMbQVWd1u77MYzJXktvZPo1uNM0
oM8DtQ2686q44+ct6dtbRBpwxCzRsGLX6obpiUH8vn6+n1mGjBz9HuRYVWuz7meOY/031imPiEn/
aIpGigemhiWmc3TXYqi/7nsICOnVBcBnuR0d3Nb9N+6FwcuUrVnm0Kv7csjX4Ag1LbgbwELokZHQ
lCCbj7At3xsX68dZ9kxaJ0e+iJf076R0aF5dCqcQS2yrsqVP6ReZ0kQLViOYXEPXufbHyrxBMT8f
M5OQq6CeqKc/MQFQifTh/ow5kuRRniU2oUFlJn8z6DuZ1EctqSqdo5MB7sRIKKla5RCKaSWhSGCD
bwnfxQHMPaRmP2Jv0xgcXWtXhkEd9GSD82AiUb2giakwxyjfOuZi4jKzwPcD8myeA+m7l6gNBizS
kkegOjjlgdBK5h4uOyAy1v+gcB4HUgXAxIvILQQ6sp3wWvqD7hzThUr2Jcb66fIgasQNfsnKJOVE
HlKR/q/s/MgVy0s4yFIUDvMDIK5z2o+h2t2eQeToXTeu0yd2fHkULQl/U7GDeh6wdht9T+UHxDXv
ne8Ty1xH4sIdAIDJkhdH7u+jOxKMEi1K4zuJQm7CXBkbAnR2123XvgVQb2s58S05vqJT7rDoSgUM
jRuL4j8skQ0IFEQf7pS0MBoAS9p+W3mnG42pGE+AT7n+84hibfKYp4DF7/vGwupFv8kVzWEY2fuZ
TRGDOj5BsCP7TUwyZDMP0eJ0xxDEvBdRsYf+OyCCU4+qDGFk8QZ0tJaPJ4zniepyQkz97bdzJCM5
VGIDocbmHhtrTag4+zUIXwXe5gBAIAIWzfJLy92G7aZTYAbppSY8pPi9KH9vuJ3lcbLkz5gr8ZMX
cB8+9Q9R3XuLZ9X1l0gAg2beTGeeQxed+BGEYHV8WnlRsK2jMqTsai59pXvcdgsak+6wMWctYP2I
N8CiRWQxjHUk7wGxE7a4FZ7I4TYGrgjPl/d0B4DSv0FIM5k62JuA3RKgJKbPyKsQTghixO9eTiH6
aSL5QH3ZqWl4dFN/x+gtu3mtyI6/q3npyIIraPeAfTu72Eo3V6t9WAzN4YJ+XRZHGW1HGAVVdCYV
xzTZ7DEeEdoE+8+yE+PpBa/hWu4g8ieFV4hG+kO1JRxmghWUM5/BSoXJtdTsdz0XzPFEGQP92NGU
ZDA7WLuc+QygoXxHR4dw6zxfRPRhAJKZxaiJ8aPs3Gaq3jPsAVqKk/KgypHxsOT1xfMPmABIETrv
mZSQwIVA/a4pz3J2jtj878EHVDGztws+4CMMwNNH+ropdF8iiN8RVEYHaPEUy65IOna4/FygkJre
1UMfAspZGTwiuGJ17xvLAYDyE1ZxUwby3rmp1ur5uOyWgHdml+yR5hflt6ErWhtABEgrf7SOsnWQ
jJOgCXeeRSpTJrY7tFZMor71FyOf9Ff1jgVjPjrhH0zMgOYtBrPR51vqlZH5LWP3dW1zUhyqaQlR
dQcXMWXLbWZBXfd/wasJBSxGHUDPH+gIdtVrmPO66y9uAvWyDADIawlQNeXZE4t9jKazk7ONi6b5
XTPWQU2eIE6nY3v6QWQVvGn/upwT02Qeb1A3Kjskzl9Fj+RMuu9U9C6uCJgxN60yus0siwbAspFy
lSabx15GqtqPMdcR+HzBIJzpVnkj6vhCQjAdBlG6cw2nut4F8tV6fhP/VDc9cjzElw5JDS4lF6ry
cPmOStEggEV6zVt9h83uA108GPnV0W4nw4izZw0LY91oKY7IlW9DdSLe5J2AJ1kxWOTemeCHpYTB
9lEuoSTmnvR6ecyjKHHhBn9fCghe/i/kRcB+fsCNQ3ZZ7SQ9zCSeN5gRLSWkNd+ym3VFZbcEuJf/
rKY4HcWrqrMkg5ROy8ISpN6jZsJ3vB4djrgv9LaoMTx0qYIcRtDdJ9pzKsv2YbnlTgtt4kl7ajHi
SoeaWrIOYPovqVNzRooflbH3Z7UQ2AkJBD2ZKCsHFYm8tXqdpiElDkHMhfxpBrP1OE4ciFfd7CsC
vtf5hwzKv/D/0/nSfgInuBVy/52cOz85ZvXrHHZH++7cRJ0c6+SElzl81FwFH+tInNjmhc040kin
kmO1kUPJQYjGitJ8ItVu5srPMxpKquSYKP1BEyaINR2MSmj29Z2VNcNnUR78fJZKA/Z6uwx77ZIw
+YXJie61YoIt4IgkVtYjFXcM9j4G2gk3cF/1JoT5VBoWXSqrosbTrDgqr08FC71Or3Ig1+y+8tjX
u5gXGRVOwIp97nAA25syJcLRIIfz2VqOa5iRgyvEA/NuMd8Iour5/IcZLppvo8AJfGyYTQ4P9cSo
APc6upaE8P2f50oU71UpliQzlu52voJmBGd4v1rot09PZ79bHE2Bj2rAxDgJ/sFjARRm/fEEYxM/
zTagCCUkUVgvCp3yDNLjavpGMisT6wQb3HV6tdKSWxHU848WX4tDUQ3HMXuCDg/bnmCXMS+tcBiA
V71uBJ4yb3xuDd8krOe8/H/Ya6RQoOnNtb++0yTKBZ4e1bUoOD+MPeD4EM7im3aR0VZCH1r1Gmfy
ihAooyZpyrBizabmnfATDsXKaJKjiEdfzillH8A/pIVZCDDLa7H8nECbi70dGtHXwRNWg7TYHbeC
9yKm0BpTO7utvwaWu6gFEk0ZqrzsY5FDGqp/0Ali/yR3nbT502J+E9iCeL0mQ1qM7hyPMWwvPD1W
IRqPA7S/g+tU3Pvabdzz6jCDrnoVeUVO2S8jHUvWxUAenL0zBYmeCaAvcRO35T8ryTvP9hZBicVD
jNUFAFgy6yLwQ6vLwEQusyQdYIoDtxVQAmTSqF9MvGGOAZmQMVbGcdRoisgtnQ5/PwFByeTY3Xp7
OqlKC21Apuzoa8h6U/AgYMczg6+UIBkpDxidpLYNYYOdZpD7fqKDoUblSyKwkl3oR7CM3H/3S7Y5
TYkAHwZFWgW6vZPgUd5m3TE3q3S4zGXnXqVqKMy9HgcMxJXI+YgfOyRvzQT7l2ekt9Su31CJ36Mw
uRNQ0xtO1dAerKR6ouNcy9+jABWf83n/APANxIDA4WHlZ0+7U9hTspeGxe7xlqt3ygXGpItMmIBj
F/FtLNPfYELqUb7fkWs7922UWTSTjIQ1lKhTKtdvuYXD9XWMkvNLGHfJumfUjTWrZW1qO9XbRo61
oY/38brwEGZyINEMK09l2OzpLxP2sEsW53pnpMS1U9TmYwBv6iDJ7lihd2vsKmjF3v9E88YYSmmo
KxFoJqUyo1C4KglnpwVU9T7WVaC2fUf8fP8mPNytvyjScvpefmud+upWPWy2PUv1YTtiE2CBgCF/
9dZyfTFPzpI0h9AsO88hh+r+GT78z95zIxgaPZvJJXHOtMEcAQF5EZ7CCdv28DKfFrgVUpcqdji0
ck71z8X/S2jqgvsez22VrYX5cdgCWxXvrbrJT8TLTyI9q1JrcEBNvakoCO6UOAzzeZLBhMKlb+V3
k9kKXYe/by+2Buu2ivry1Y22dv+QxyqKPa4o3tXtcERkqlv2C0x3twMpZ0U7zROls4wwjPJIVKm4
0WrO47P5TM1eULWCOkquEIkHzPGWIv03jq4SlPhYQPIye9rl/msbCqGo/5anHI8N+V03E+eVF50+
dG7tKeKcezKuEOuN8QN6qxkbMWg+/K5/IU92/J3jtQyvKG07wXy+Z+FKH9iFYxSRjZ0eCGL913Sq
dBeBDiAApUf903kr98or6L0tZ2woFxFV+CNFCIUcv6xQ7e/FVkWz3ddHkisUQlUOVkFqYwQZovI+
Zw4DOObaFEBXdN3qgVt1/qwO+awhlkCQiks90TSckQvq9Y5x6Coi3Oeufx8tqW4Dr9QrBJpccoTL
XX6EXG4fL+fKnivZC4aOxlXm01UcgZsIOIXptjB6VwiY8oV0NO0J0OZEzRWy00CY+ekbSuhJZpzu
oBNHR+xWembuHciYCfu/ILfq1BVUX2DGUrZ5BWaBy2gCpgZvGWSpHWC9rNs5KAtH+Y1ZfsRxmigd
/AcvHFAjyYA43A/ZyzBU3hrDEOzKjLek/oi2DtVRWZ/aP4cPr3Antu8qF33GwAPJFhMlxpcWT86J
fs3gYuYFqXsrtZJMoSHRcizPyY6ri5FWxG4TrHTqjIs/3dsU35//auAsXYS5OKh4Cd91chnUGhgq
XHQR94Ww9DVHUNuxjI4h+oadaeTtwjSF9SAu6MWjd1sgtU3+r9fCbxvMY2Cs5flPVDtYA0zv5esp
6y9uSfbfqdLz4XDfhKhQTzVaWJOz58NYSucTin3F3UwqfYzd0OGqHiuWslbdzG1jaI+B3aly+AAe
iTldsgua4PudsCKNVeO/NMpeqU5aCJ+WWdf0usrRdIMTDNPAE0hAsHZHWl0EaqzRwP3/dnBAmUdk
oBZRviPMwv4Q/m2gPXuudimAQj/KGKOfky7WNAUSpzn90BRjkJcWOS6KQf/43Bhj3Sivz9wxos/9
Sn/ROI+itXm65hiDRCT+G0ndUGlGiyh8VuYtjd5MkX5ABjtA9h2t/Yv4I5lwyoFIUQCuEFBRDAVA
f+DmXmq7lB+i9XOYOlNLlwJP1pj7aASGq3IgKsw2zys5clivUYomyj460vb1hbJjhZ+TodE7Bu4l
IGtOJ4Q0XiXsVSHGx/6to8MaQcOlktEP39/EiVQeYX3yuWsCRNxSo0GGAZRnEh4A5A5Kg0ASAxUZ
t40CO2XEXnMRDTykmTphRE4PxrKGOR2a90IsxjBWtR3TTH4gd8sNuKMt8+N2xSPjaV8t34eYR7CD
0XMI9EhWr5zL2lxAUWyOX7nN5F1oqOHbBkTRe8BvXeeFFiIhLDYdtkZlOp00vYJKbK1n5VXlYZ2F
c62ec8r+Q0qphqbWVj0OsF9oy8k2eNutoEJGYR6GAtIYg3iFJEjvVq1aH7YVkISiWiNYPOiX+7/A
kNcmFkPkEz0Gxqh0UP2RFS1Yo8ksyaMB3kFIteu50sbFK0LrQg0IUNS/58BsbvdI7Nzs15uFldIo
6deyRbLCaNPZIXldz5i8TB4/zJFeybw7oZFgs3I9MGe2qrQY4zAxujbXDGi5N/Dmt5AGW27vEjUG
Hajwb0/avwXYZrdoCZPu8FP4mjb0V977hUP12ESjwAHLMT8L3ATRC/v6r8bkh8+l/oT1p9XrMT7n
5Tc/cvgRtjIkAUzZCWRtbOWAZ6NVG2RMntaIe+NSgtLdzy4Jdaq3RWxR/Evc2m8DOGgwff1t5Dq7
gcBKYDz99gNBhONxj7Kz72wD1eefpbAWycP13lakjwrRDMJQUX4DMkAzWd2i95/r4KfxZoiTxBLW
FznhUNsNmtU4gXiIcWWrY38B9H7FxT/mRwlxpPUX5dhf+2RVbyxGAqW4/ln4MLVg4E3RBh9SIW0m
mv9xaavxqoXOaGPbyZHaxnNSAUFq/rbJB3PMzWEToAqguMNv8md1Gxi88+q39HzGd1qZ1Ed6F/9i
m0YiRUdDhYpmRrWybbGuKiP4O4d7KfhL+PhdmS4wmOgqorf22EsHo6ZdtrcF5Y1BXMIoMGtcD0kT
wMtSy23jEVw1EybhKdQbIXocSPBdumUMfAopmNgIckxKivDPe4wCHwNTE48DXMa3VMKUsNRK7a5M
XG53p1IzX8MMv/ViTN8lR9Js5T/A8KZ1gQGA4bkv5gWxcMgSwKzdYsvnY60m3HUu9Pfx8h34FO1G
aFNHznNi+sp73tLC/7Qvqn02YX3r2GLtZWIa09+jlg51K5rOagvGDL8PDAq07BSpqSCPCihRnEoY
GbQhgJoousMVScupOBS2QWOd4ZNSLQPV01QN/0e0o7QI8qe8hj3dZ9bJ34N+bM+/TP3AAsb65fwH
RkUMXgwlf7rhy+8dq/8uTOaXp05uUOoQxSgiqQrpY6byqBKzXfMfCL9nbSF4KXmzmnEm1A6p9R2p
ZazriC18dhkngZLDqpEOV7fpnDxEB9ghI/GYXo6wIlattcZdWjXGetzIQrAup7K6cG24XNHdTWlC
+jgla6nRGqaLxG/m+GRPP2BCWjsWJ6tDQ1uHiGOxN/w8Z/W/a7tL/FqfsusRvy+4C63rfHLCJ3VG
21LuaMjVSKYTzQYCT67+H6ajgWFIY2FWrki1UOIWpS3MfuYvAFCb66Jq8DhS/gRsFNeeiTDqI/A4
Np773BWagAQ0WqwdMcYpctwibqG/ptVluEllpOMeQ+0nVmIzT9oH9zZhqpAr35EF/Sn+jDeh7yCy
CMQf9p1bXIysKO/5w80HpiBuQa+ERwUSjDcWO/PrpJP845md/lazqGCPbRokR//Pow/AWngwehX6
uuZRsYl5VefzWE7lZpmBmnk3ygCpeJ6uQTO1QdqRZLFrSIHtUAUV6Up0WExrA4hDKpqzmkwPrJxd
Z5Wcnlnvu6BdYdKUeQcDTJWUQF+yzPtvLDuwsNw14drLk3MmahPCDiIza+oWoEgItdtDgsPaVKco
MWNxh0ZR8iqVfDbT4MJGauDTJmVZG1ixahm0I0k1dv2RByagNt9FQ0TM73yC5tO480mMZkNPZ+LX
Gbnc6wq/+w2byvVOUHe6ux9l1wksUlv++kIxHN68RuIJsiJ0BQcjSrqJ19MjAXYk9IldCtLBTzSM
pNYb4CLWKbMAUFz++AzNzqew/geBmBHaUYEnPvKu5NmsjbdX33x3j1l7aN4qt85KqwskyzCoHQ3n
0RIEMJ54jUu9ou2nkKVd1IojyBFr31ZSvbtZt+n1piX/KuJN7vQov3rRUrr/DSYsXORbeSKEa4j3
BVD5o2du/d8VcO99I3lqDL9sxqALF+DZ8/UDJPDmn1W8z2UL3zyydM6Lz2TQacYOt/DOagxem9eJ
062BYk29XTewo6rdi93/poxXboooXKFji016Tq+oMGWg/Bdc/Rqp0EmC+EQ0uoM1kVIFbrl7zy08
T/FPdDfa0vl2/S4LkiMZ4B3Fu8HhuStyScdeatawytAoy1DmgapJ/t/EHLFfFJZ5irbHg934cbso
F1dKb/Z9b9iwzCemUw6RUNBj9QPuya1M89ONog9JY7Q0xGY/YGK0e3S6YswjMQW6XRTay7xmPQmo
Wji4EBrVctY47C5aiXQI97dyOBgojE/8u4DWj0A90EKcYreCtWOSSctsZZ4x7wxf9y56ZY3i6Wug
lgxjwtKbp34AjlskadnsgaAiAMi7SaPXZM2rV+QxhznmnRaOwxGZtHgxUK26cpV2BgKC2+7skV27
4VWFOK1HWDM9OvfUnyB1B5YDwnpSk5n8tv1rTU1ExE9XsDn2oLiB1+ZyMIEeDYpbIZTxXXnrnmdg
0omnngcv6F8pZuqrH43477pKrbDSNdc9aI5XIdasir1HOckaiEh3LZ+Xx9T5q68mTHG4pxXO1dFA
rM3KBd0LWEd+tWPpMwHu4q+6btsWqCNeUHBnrcywrki8p6XQpuVXDOoSvhxaUKANwOcDhI2DgQFQ
c/StsjID01vx99/3smYcQ3nMTf7/Kd4/CjgzPyXhr1qBG9kvqQ8A1+oQVUmsFe8nYcCoqG0tbOC4
An8R7c2iSgQTyICL3TjZyZqLN4qM19KCd7VZo1CjKNBOrCej2+hFZVbwSRmCKi6sxdsX/9phQe+S
ScmsWPWjMpEmiJNkK8OkRtyc82xc2jlFKW3ZNfy5yngiZ5yJq/Oep+e2VixTTwHaYG4ZBOuGUOJE
bAqOXuDWPVsBj20pqPdAnHkAi3JdYopWR27gbZwedkQ6JHs3PwbHT4GjcJs0XarvbrE94ZRLjgIm
Co8qKpqTQiO43LjqkZUFK5sMBYKUoSUKSv+cyq86H7luM0Iwfu4bOIVJ1pW43F4uOTVvFfjsW3yN
3A+U/lb4YMJKb+j9WHZdnbdAHYZa51CMoR+D77weyJ4uIeeudYK28cwyLxtWSUZWtCV/anpiMqBu
JLAkIH4tR0rtP4UwcL7uE969dweLi8D3P6vYt7W7Gv8DB5m1XYhfHX9BACnmxMeHmz+Kw76qYTPq
DHkjNTo4Qs5pcplov0VkYups90TexBZxkrFqWwRA4UlBzeyioZkKP6OPJmrRkgDgokqrN/reipTS
gNRss/AIAWrstJawSaV6FcsGtEgh0oZiHknkNBGo8KJwyLMPioGlXrYnjOduqZbExcxu1uV05/WI
ABfSIoyS5As2ZH5hP6oKEY5mdruqwgnCumeNzkEepMK0UE6PH/zAt7QkW4+9E5YrKN2KDXbbZYK8
Gr9hcZ6UMbbTjAl9UV93Fat70ltUkvWOLfK1gkQ/67l5WnatWdLr7cNtylXXrItc7Stko8gffGtM
9UP/Rx6A6PiEDfe8aLLo2LFnZEme+EBQDKq7sjaVHdalaCtQJ3uHfBPPbMe4q6CmrlsXyP6DNJMw
vgyenZwcJpJzVIrAjCz6rJJAFeUdBm//bdk0oZmoYg+TVAUISwCkOJOPR88xVHroJHuvjGSQ4zl2
OT9Vj4P+o5o/XoJ8xFQ1d1HzizC890lK2jRdyEgD7oyufIsuseLJxpmExtp3b/98evW15076NDk7
LJAhcvBWh/dHPNBAWT6iVkGX6C6p2A4A4x4FcPTJo3P5ytzIHV9kkiWz17HrU3Z1ipZNZA5W6Wym
j9qwCbl3/z8zRZEXoAE04xrReF71McOwuFLZBu0icHEnTXXE0phFTFQa9ODXiFkEBnnEURmPouep
BcVeCrEI+jLoYwqcNEQtVEetFxQbzjegYAII5lWlKuEsfkNTbyAzg6b68pIFmXCoTWEI1A7r5gmS
U83h8Np5Cu+b3ClXjg8djlLzEccl1bwPFsYZEi24Fsuf6kEObnbEtAyl0yKoa0hv4L6QLcSrdaKm
TCZjhyg8PNacg2ZHWh2Y0VyI8g4RUNLx2M1Yo7E2XDez4JbBLqLs6hB5e4rIyKpEj9gTGIVi4KyO
1vgx5t8omMN52WXmHQlq2rBTPQHILAce9zsamu34XUDlVH15Gk5SczIpeIYTlC7aIvNWi3svbzoh
dC9vnRkmI+y2kNZCH2/GBgm3PzBirKT2nadzsK6aaOJZxTpbhOPSpf/y2eb+S71XvxOWAoXnXLKQ
3Qw75DrtJnjkSEqo0RnBb0AdbAX0sy6ZO/1ANI0nWrKqrHSNhvK77aYLrRHQ7q+F6P7/n51/iEpO
WeFkpf/RzTRnhVum3oMa5f+TzjPzqG8Hu+Hnb/K6TOOoR6lZxlgEH6HrErNBO3Hg9YRhq2blzS6l
+jiMDkfEQ2MG6HfEoPDA2j4NbUDE4cg5aYRjvhXjK8HHK2+/w55WfibBENK5uO00rhOrvBSjGfkT
ke8CJ+vBzfL1VgKsF9yKl/30HP3ncRRR/k9K72E/h9b/O4Ca524EnrlB2BISL1VlmqGblj5pUISL
BLM8jknmH79lAL8k9ei/Ey4XgbWxqDDI9RoRZL7b4qSVjc3MNlHqvU8MN5VXIGDJEQWpNSxYb/PD
N36tB845uAYbbBQr/MoytNW/FdLXV39hBPh/6WSN71bMRiHJLDUqR8FZax8/lVTA9AoZnl5UObuX
H+g/sk88vJ4BXMyg4//bTO98dQYKn5N1Rd0NXmjicdRTDOO0DIukg3vvuZ3YYIpUppgP5wb9XH7k
FoGkCoUU2lX/nz4xF7+TaEblExknmwcZ+f+ha4YfCoBqHhwZAxl2I0DjjOy5fu2IQf1VhBYSy/5i
OkBcOom+BMs0r/d13f1oU694N0XT6MMVc59KBVlOcDKknHpDVQIdm3LE50aCOcCwfg4mrVM/WLgr
ifamtTzrOw00+7IkM8CTLnRo/SsEhXM+OpzB6xg8uBrd/4nj5eRpYVGBoyI/J2IsD3l4AzVzLDc4
oGKiDOFilmEVfi9udI864qCbT6F7hdvqoKBgzfJqwfoLIM5Kktgqwu8ZGnhkRBJxmWNwvQDhMz21
8GfjUkDbpkIw3kW82+VVEwrmYgr6lobQ27r1jOeXA8Vs6/kONVMeEj5j3nlT7AVEtK6W4Y6ylHJ4
KDK5FAtmhfz9PfvbCkxdN0Jr7rT9jhTn/oHrtVJjj2H+KcPO/sX4K8cQwVe4RWbyV1kwRtZqMoOP
8GxqTrLmv1PILxpfje7shpo81cgLrix971C/8vzaR4KrA5zBsgz8m0UYPgK6VidNDdtYYFpSH3gQ
ox6uRNhUXefoHaZlhIaVGtFbZreb1L3At+e3VzDJNbWHvEWZsIBjNkJ/J1Hh0eqYW12bYmyFhl3z
9hmZiInwqV7sZp/lKrh8/89PHcvvLKxNR5Mz2ANRlC+vhtAtsvHU9vrp7hxpMXgdBDvdh8B9cWJd
8O28CvEZTY+debfM4B2R39IamqSdPT+EBRD1WQbDhK39K7NEZbx5HR3CR8lKg8UFptpJUAi2kZTX
VS7AfoAAHqCEE1j+z0KOKmNycoVSsxEfmXc9c1IS2J5S0SLFsZQhDsdMn4SbqZfpkdK7lELT3e28
j4Jmnim2vGEHgCcb+3FyPudQMdLgdNXn3MbufVzv8uqs8lzmN4C1DX85znAUaMQUWZ8h+k7c++yP
ZxW1QLvtVss/Fn0kPqfwIl1oelN++wFY5/fZ7E7ZTp+aGul3gsrQLA6LCaspMZhpQNSrhcjxNWTT
ZTq7Qde+dkhj5T/LdDZGlMH0OA3GJDUiWxeHJXA5L/o+qUJSbYKJv5jDFQm7yO+fe7gtwcicM3oi
yuDMgVhPOymyA49Ytvv5DWDUGDbvJ0yaF9smpugTsnlrL4bgIEZdcucUHUrafNVerG2fI9C8BaBW
tQgad9l71VqAfvHorgkdoR4q/kWq0HQ2wtWHySYMmZwg3JhtrDLJf2fLcv9JehVP6RXKfDI0EESz
ctZSXJPLoGmYrYgzxcqb6HHwnELoipVq6zQH71W0aEEHiso9dBq5E+2pObJIzTsnt+VXv+mBOme/
e8xHJ9s1j0TrqVrVcVz2gGVKwL/95FpVBYXKmJ/Q8c5u+c2BqUJ0OcblRxP6zrBDIBljO+eeG2uq
ZeHSitTIjO98rl9tN8L4Si0AZCVK0wElUoZcI6a+d12WXErnh/WH5eUh1a/aeJHVZXJKbzCBn3+h
k7EBBvjQqg5r90vfxwKGni+tao9ySn/aLQ+Ahcr+xYkbXOP0ankPrt+R4uuzYC37IgpL9OK4D7ng
03Ap53RYsJy/OfF5kBDqBa8Bd+1l+AMzNO8eM4jQwFambn6ehS9AJDaczH49r0qn2odMaEVIOr6E
9aOO3zhjzbLImL040fL4a3eSzU+R4xit1ERyAxeKDkZd+QouNrr/fYV6OUmN5SjmxxY+K/4vDojv
oAPvhDbRu751oxxmfugCJx/q0mN/Xa5+qtbZ/EvUjYS/VKQRKnQ6Zi1oxs78NjEgn3ct87jdZ/LH
WwQZJqPZlELccXhkNIBPMTQUxfYdqJrk9zxXIwe7GzEqyOTLqgC05oQiDrvx5+KCDhgjaZCp1mBq
s0pOSMgkRjlG68GW7+DgBpjycp/WaTlCMZraIIxws8MafqElQRUEZ2UI489EmMOcCPlqvk24z+gO
8rHq+wHxX/7IQAvc3e7qhZPnAdcUuZGLgHS+keitbivkV8DQEvq0Bvayt2/oE3TbEaVDDrAe6GlU
l49mJgUD9FRhG8MeEJzL9TEcSrY+/dBOalThatZvBucIzr7Bn5xFRw1uKM6fO65DMFGCTUHGVHop
k8GeCENrtqRumbZNlD4VaGiiq0TB6+EblyF0sV7xO/uOMngkf74DlxyK9tEK7xkmO/zapnVx2nYB
+73b+t8U1m2E+V9QDewSbx1PJE8ssYmawbzMovFjUHgj1S7OHS8VA8W/Hd9/9PwEq+dvHcam45WW
2eUF8SUqJPqW5DwKmlEDeirUG/bCtm3CNRCANR+AYY00RpK/aQl9/VicBwHkD0SBor4l0DU2D6RX
aSZNNXBR5+BrWtKZI4fn702IkxU0EffEL7CgDOw9qxh7WCvHiABjWs4gfSD7TdZfBdfOGorPgJRY
XC6jD4CiFEkhQG5LlT/nGVzJ9Y3okpjngv/5nGx+QQDOky6/AI4f0YvXokTlTT+ciyHXvdScdn1j
NFJMmLoEu92ySbtGBH+in6K5xahtSfoJk5X3Ukqrohr0zBZ+9CIOdVzpH5WD5JIgLUX4TxnmAUx8
EKluwme+Ar06V9fSxxHMjy28FDbtXQdACpl4YVutid0gxI7NHJ9LG8kxg+W0vjBrlWtGHBg3+MlW
7/oVx7Q1QTlyBA/bvsa9Fi2H6D19jW3C0KuzXmPDFP7/NzHXShUhTkaLncQ+JWA9ZFseFi30p/ws
8ZKTLdW685WjaJnY+jIQ6XWndUjYwnKr3XVirbWzbyOJwv78ZDqEAE6DGIhAe7PlvglO+mGemRkL
BmfKTRHnTakmHjYfh24i3FVyxbO0t1yu6I9QZP35hdSV02rucBLf7CBMbk/FUVWP3dkqnCyR2yk7
6tS4C/7VuztqiKgefcfg2jQFQ2rqR4HCV2L5AzieGdQUDxGapgdVLU71PWsbj35/Nk+dsmbSurB+
QdRbc6bk7NxifRGlkbS7sL3I5uw/Z59GpELpD64qcIwCGPQjOqRc6nlKbWt6YcEm9IxVBb/Bp23M
AV2qd/DEz/3ztE3DFnvYyylG4cEahbIUPN4E1s1UTzgzk13fNepPGvOT5xsMfe1WDRPJsEFh5f3O
zLvHMXYze242IhX/hOvkmbmO5VG4k/ORzctZHV2BG7CuY2gvD3YtoxkrHkdZWX6LuT+Mnu/9dgx9
OjHV8tVbUZ9uREgBfFYXnVymCySNWIrYy58j4JZ0EAHc+WHctSkdggVEq246AXp6q/Or6OzWEhmC
2DSPzECls+V8BnMTu6x9XLFdYW9AR2b0fVbFDBfMDLgZNAzitfKWVl6aZTjYcelrxnyh4fkWr2DB
xQIcnublNk79tzvbZFrZunjOOJMKkUdztETu6huaxTu5jPj8B83+MFaqxfWklCuuF/OqrpQEcPE2
nDPqp3scwWvRGzlR9CDGQTDXIKJp7DnzZ+UCfZRCCeRd41UBLy9QtPrJlN56u/I4J2Em9aHEuJaZ
SfwoAdAjJYLeE0KwrIHSP1G94k8KBID6fNzb6mU5K9PYWOPwJADLLpZiIZ4Tp1FE4C1ES6A5mone
UEskg6ujA0ud3cT80Pjy0T7pGl1tyA4vwuSrj8Yl0U67rOZcChdcSwl8NmCWaV1f1VkVSu3JxUmK
C1w9tYwdEcFQO0mxWtGlGyjbIur2MpxUOkZrPFvEo430IqVmkxf9suzYkQ+M+Z605bk3M976f/X8
Xj5olmdinRtoTz9885BZAE58alpHFfMY/l9rOGjLOO42buqQ5a9H0Qrutmrhxk3OiF7iW0ZlMcLZ
xHzHHZzPCfx9sod+UD+832pvLGfOZSPRPsBF+ieGQpmtkTr+yRB0pD/97+opfCynqALdKM5NG6aI
K6+jfw34pwuF5llo87CdNn+N6mZy7oxMQimcQfUvKN4XXRcxetEEwbvLYJjyTkKzepx0UL0WTjuI
fhe4bH+r8h3A8vSp8mmd5Qnfqvezu6m+4SYoSjE3EU1L5YZXyeV/sdJF1zswcPnug0M2p/ip9H8M
wR3jg2fC6ZRblP2Zvb67XO838gua1A5FdBNPosnjjKj7Vqg01zTxWoIAd1MjA/s1/u9HbntnomoF
cxPquJBAkKyueHTiGGDqIQID/qJqJkmad1MC+ZKi7vc2TZY9aZdT4iVkIqc0kLoG1c93IKHFLBkC
XEWIk59rqHfxKIBpDAcl2Mg7bL4QNWrgOd5p/wChbbNvdsHVJ1SmwKr/Gr/uoaDtlSu/+mQNWKoT
kB2uGVWhm+DhbZk3G3nVX6YEs9qweB3WK/y5dt0eZFZbMqPEzufpthmhJpjMEQbdsEMjAg7k3Z9h
ZEZ9okZWqZrpxtj3LHqGn1nbrWxSncRiiqaMFC5fBpWNZwqu0MpUwRdBrERlm9VnyJ5KVVe1Q982
xuFO10BWoZJCSX8MwSm8+40wYTSsZ98RvUeZgA5e4otqiWkhoXX+dwHfe5Q2wIWfWTD9+EPTPq0D
1IKf7+RNyc5DdSQkpz68CY5T0nudULbaS08rfG1zhz53RhMNB5WLkav2zI2Z0CmeqHvYhrgpQQ8s
LNzSDKfYFgcYRK/ymcD30zuXWrRtSRTgaizamo/eFVKdGyPNOBRr4lm0i7S6N065uWbD4H288A2W
eeStYXVYlxq7a8hgAmZl70brGmGXQHjiEqW5OVzwdSL7uuh3RQM9+5j7If/3goRaA27Ye7ws6iur
RPqmzYYvZuTudEGnbLIgn3FJLaw/mJGaFWRNwbnpTNndTPT7l9mKn8Ub+erD0zA5NyuGUmKjCEFP
hM7zsyGnMDrgW4sYT2mlq2XiLQc3Tfwgd9HaeuswVrwr7gp+LJQOfr8NQqGIhLyDbxSXu7A76a9j
t8LzY4I9cFh9GR7vebAy1tXnU+Zbg5BG1ZJ4HlwzY55amja0ZlueIYmHG9jAnZqRBQebQvGPOvO7
AKJG4/bKxI9hrd1ZXfq5TZoPdak9sooZflukLcComJ3+wbkkRthkrixT8gXsFd5/k6xRzQ+HLk5L
yPJ77lLoWPN+68eNJN5uUh8z59DGhBQPiNQn/Qh7kouUFBPkpuRp6YF1nWQZ3U7pGGZKrCuI7i/P
bNItnwKZOuD3zpRZISwoQV5KU46rZtFXybmthn+IAcNSbXQwlRtmcRqa2WxkUfECLjxI+6w1TkHD
+tzHg51HWIkag2/7euvSZuuFqR9hJaM8PffcChcSpWjQ6nnCjTezJ20edNtnf4M2iAYtHPLU33y3
Eqp8v1y0VucDtblRijog8gg0LNwIyz1j6rd8vDGpNiaHpo1xSxrrGLg9GflQlQ2UAH8aiRur8EfH
9wjVdbAD7jeR5Ro2UCfRB+nMTWmfMa6ExWFvBa6bkYsoyGONcNH0KE6qbzTwIFaBfxisZXnJ1jOP
1VqL75/5G4C5pdbeKt7QLtZpsayrsrjtZM3I9w6IIuWhdVp0vgZtSxAsgecgrGxgftWwMf/XcfOC
dxr/Kn3zPvVOCUGUIXm51qFrXTC9qh4n9Uqxu+i7bNi+geJLA367yR8UVNRcfIaoePtfoY2HcWmj
PAuAT7zK5ekKIbFFoeIRI5y73CvbleOzGoaXlAyp3h4zZXE0SmlbtbunSjD6NAkkHj0AAOHtXSMK
pgXSzpyp2jpfsgqeFFXN6nGx5ZflVIoyCC1Q6G41JdpLbr9dvtkeA0Lg5Pb0bb5Ps95A5+BgXBZV
jbOzwFNsrgC88jVta6owFxxgY0tAkVDjfp/Wtjs4jWmhUiMJ1OhcfXPiIZFH7ULLXAF0XB+1pAVh
YO81hdYi/8NdKYefc3fgfqBBGwrcp34XJCyMIO2RWJg/t9K50BWV2p82ztzn02VjGRRsCSl1k3fW
918tt5N9eWJ7aNDx+IMJO9zOFUdWHae1R6afElzqcuWb9t/nV2/InIaOrYxhuuAtHWoKu+I4u8p8
ztfs63W5fLhC9GtlEIstIk2l5FlWFJBIMFyYgdB9VaPoiXLELaEnQ0fw1Hz1bLmuq+KakavlNsPG
58ibVqOSlDty3J8jE1owCR//QZ655ogvu8edbNwE2RsKYnYidILpnnfJ70Rx4Xy0VMDcnFCS+4+w
cyQl837LoFR0H2c2aHG+TyntMxZ+BQVz/kyoFaJ6o/ZhczVMp9JnLCfAjypnQInGah8hO9GHrW/2
MZEX9s7ilUC9kka8Ptuw/vlLm+Ccf/Lpt5XMJ6Lfl2LRhRCH4ETvxn/bMuJNhUsrSFGkA+GKPLjK
Ot34X6QarjeFmtIIucED9BXXRuuSPhm2bJb2NxrNRrJOpqt4V6Rgdj3AGMjmbCXjoN1IfPf31YYb
4CMWCu4Ob1czsndw29B8z0MXRHcgJkqD4VcrCQKR6y3+OUm2V6ZW5BenQZUCD9712aENoeQjNYi3
oLlE1GkSNe575wHNgy+A/e9VcTTgJxvm1CgrDSjyVMBBTtCCm34K62EI7fMIUtCdUrT+gtegWdZw
h0Rdy/rs56niXez7BldTMKbzPtKOk7i9nkE+hayflhf8h/bFt8RYiTBCinO9eKlrwVoKVvQajoZs
IthOTc8BmkV9Xo0cwxc3S4fnugkRqUMNODbgkdbEp/Zy20WgJP/SGnXtJrMfX0961wUVqUFiVp9b
6efLPhVdeQevRnki5EVyFbGD0VAEfqYes1mq05RUfTUXG1QErDUpuvxPvmLnL+YWYsCmlvv61flE
vGnPTrIi8fKHstI/h1iufAFPZALXrkSz5w07PX5L3jcxAnPdq8TXe1Q/JeKVGUmRuP9jmAd2/9lV
2JZwA/70vgfOjz5eilytAAzzcCI/xyAvldue1GPImtbpcMuT5McDrZGqXquA+gchUN4c7y+bABbT
0l16GM/59NGkaglE2MlzWK1q1dBJKDw4S0qQPzG0lYtAh3a/aBXb+7t2yLAPDUeXOFLXlslPQzyQ
R7spU4yfOTT5C1J4+LHrN35+fhLWKGDSVj4hC5eOFnjjpr4c/JNayt/672qcueLEagXhtWqlUGZ4
99h/nNGwzwFmsmyiYO6FOlstX55JsDbOnJ0zxXUAgd1uwtRFNqDc/MDPtSJLk+8KS4Rv6y61jBtZ
QPiMQigedAEpKO2t7jDorc9v6si1N1RxkWHlMMorn6TBt4nzJQK5GbiBNUD2/2ujOO9h8MkR3HDD
B6GusxrKv1uYNnwbsN9KtOUTX80udo2iMpSUPxH4r9hH0Jxa4XfL0DAFHfsIBZMoC0x8QTRgT0iy
itD7pME8E8Tefl9GfrJvox+aDmqey25GVgUh3zpvh3PVK7Bc1f7XyM1uPz6S6ISWOAy8GZzCx2Sc
aTtV0BQIIgzbppBdh1bH09+dgQaATyOulvAZDbXxWH4ckR4u+e87itD/KEsuZhOn2QZomaHh85Bo
j3ewmexr2AqjbifNYoBed1SHUt6LPvOYPX3ox8VhSGHwghcLkGzp4BSkXmIZ+Ef7WehFQngL6XAn
gPnajSZhSZ3XlLzzNeDIE9g/koUIka1f3YA4NOViWl5P6J3BelKDeO5FREFo8EFBOLxJj3bmKFn9
a5Q+gwDvOAUj2Wa9fcfTJw2DNPe2PGuN4jcbCyKIB13qOYZaZbRsOrgmtuzhAp++TnEF2DZGKbkk
Pe9GoyhSDejl58dSnvMezNX7/wBNP7iipqOOPknAo9tkahMK+Py4A8GN+7WL8EfaBJ3XK93+E9s5
y1NyJ5YY/PZe5QtjMb0KodFz5r319Uc2zccqXUB+21ETE5k9Vesmob6AgCyCMIp3OeaG9srnWtpv
VZ8Jc+Ft/nliciuqVDCCjDCU/GX8wfx7bmcWhiBWMPEHBw1FwmZBw4bFktsNgqzw6UfQcBDO1xzq
6iq9f/g+vYNVJo8lNzVyfD7MuwhXUaVTyQd6WxKVmdl8bOiZeEkEsgIxIr48Xcn/5D/4nvkdXZkv
1Z3WKyxRX8WkWIHrNRimgDJv5RugP16jqujDwoGxnsGBOjm0dOdweJLQgKzxyWmhgSgKNKXsP9hM
XXW5UsPXf4dENiN6DejsR8ppL4aERnAuzWQEy1cXxHw6qyGSmHmWt0AoCV8SDmCwdcrgOjtEn7TO
NXmE9+1FF7LZtbjkRWk4XYbONcqQXJhblUGX8TnjnwNZrzQuLcij1iKZ2nMcH80daYCbeCeWmZzO
wCd1Us8oKWt16T2jAM41aeblQ9A5bX/otJOnPH+pMm+sZYKcx5cklHQ7Y4+xvIiWdVLZntsv9wpl
Mo1UYV6z+CibputM0OD0WjyK16lv6rn3Pq0CeqovjxR8UH2pmLBGbYHSe0zLuvQQYeSgShdSQp5C
Fk6FOkmdhTpV490ATg81ZWLqWfgjNPc2BN3GF1t6LhB8EW8iGL5x22Ta5bJlbPgsGAIErsPy1Qr+
bB7X8hfNsl6jy3DsJhc/84/jmQRIPEH24RKKDCVrzusqVO4hbZO15ZD/LrDAqcLVqeG98Nw4exI4
e52x/R50GvN5geqvECd/BgSjIiyHftTZVt6lnsLU9KusuEeo1rZC0PVRgYaUpEFTwK6TSRqQQsyq
TTc1OcWxtxDEkSHh9c+t4K/mhZwl4Yz9fL+mmdSvDVdMBmhA9bbwxkEJX/rWp/rBB+6bHJTK9P8s
bVbecGT5CIrDD+dZgNYKjlWuBu/ONAyXjangmULFmEyyuiSMojUMeHUmbRFbYwGQq+UYlPCjz57X
atlVfap8Pl1lBfFlf5pXUUAdMrBnc1exqL8NOu8wI30KXSDDH8jCr55jKa2upLGN/Rdto4E3H7VA
c/o4TrMhDlkzhixu8gvjwhEJwJxkKpp6hS3zIEADfN/4B4tZw41QUJT8vNR0zRagRSMr4IoGnPjH
qQZAwFoPrjnWZN8tfYxlQ5h01co/NKjofAIUsBQlhEyysD1tOE8vOpmZ/w5T2/XuNgk2ukgKRdYm
pkttiFEpfpx0mr0pxloDj6WvALMgIocLKMa7mcJHhmCSOo0e9SHGwZeZDxVruWFfrG32RmLLGKiN
o+XkFzPXmak7dyKtgz5vJFS7QmnpkGVpra+py85EbPPd37O7okyRCjMqusKSFz+uj8Et6D6qXh8n
4/evWLhjZTMjQ0QMpmTYxa0G29LvTtJO8GlhD9/LQXPEeqP6h9sdO4TW9hWLQcmsThUPq4QXRX3v
S9SVCmDI5NgxlBeuCrFutgX0v1w+mfs9Him7YtDDUCXwKaH0PSRBvcMOKDZ2khwMZ6JybKCTZRue
iebkRQzBzRgdQ7CbFnNSTym2Ju/OO+W7M7vOtke+cK+2BoOg9STsDSVjvXf2aVyGtfye6UeY2m48
r1vRiG4VYDq9biJV2BTm4aHbmufQgz7tgqoU66zBSrCfUxRSjXPmLyunK+svC9P+P0OR1j6vVfyo
vgKsnNWRmYCmbaaGT8VgXpfdkzr92iFCN8HXiYxybdaDTdwdKq3/4aPmSBCqnf2U9hH6T/ekui4C
iyWGV/q82QeIfzY2P6AHHpG6x7Wv/+qv1ncREEVYMWzbcJlOyoM0OH5JUga06blDPnC1iLmkqxfa
h0pm07wbo+yh7x5PP56wEmCaoeNeny0LLIwZqvL+9V2e6a/9MEMbzYaK9/iQwB5llhnXopLThzEZ
a+DvFqEMLUlaSwIZZ5yi7SL66TEyXz3KTbdK7R2LKrG71oQBNtDKpUkhZ4U1EKNFIBM/JIsVLCl7
Havy7OpKWNUJNUXZKe+Bfe4P8aYVuG1lQcy2q9PQWE4LpE+KZHG7rarB8qbxSmJWDPGigQFdoau6
pLQgQgfB93YzvFogE2Rh7xZ8+Z/fR7oKO0FTWJ8nT2NY9loQtauLuY2x2YBYXNb/NOsVWebqz+9N
ZM65VV82NyChnkN+gaqWVA2InRrw8iEr9KazZjwREbG7NJ/aFvbE9gjvkzZa/2y0BdUh35j1CkxG
tAUrpK2ebiE3cy9VRqredvEqqetQ41sHhnDfov/+RLtRJVSMn5q7myUegQbiUN1qAfmcRq6vOtxZ
lvfhV4NmDp6s2HT23za2/D+4bzrjfROcEZQRfT5gq8niEKCn/S3nBwvYKTBxh0C5peWuzJm9XDi3
LBzUv23GBeQyz1UnNf9EO7/0ETAA8YkPsdzSw/dI/fCzpIYLRdf7yeUs1G8XNrDc7vjGEJyPqYXW
gk+bC4zCalMoAsTy+zMKTufkGydAz8aLbqQvBTuFuvlLAnLaAZqFU0vsTKB94zvYQVCz6AsjcHgS
FbtWqc4XvkWMEOWvczaZYCgjGNW7rD5W4oLIvuQRWCsfPwjTCuQB4TzQcZgZK+rHWKDaRxrz/64J
NiWqpDOdn3vyOtWnMl3M1/9zJSMW7sxy/6n7+IGJI4+dnd2bXPUMd0RmIFiPkJVBxkYfgrd/aHFy
HawSFLsuU/PKvDEAizlMWZZwy4i++uv7fwhrUV7Xc7IldyPlDpGsYQxd8V2frBdcTpWAiTkX9BH9
+t9cP+qRVxqES7tZ+xkOyqlMooU+MGFvo0jEwN/dLqRAc4ppKPoXPdbt+oTXvai0H9HNzihPRlAt
m7GmEdDF6FMnV8FUOOAP2enA6BxSVvzyISxd21pJcefTXJfvnAwqkmRugOw0MV6nt0y9m30gPqqe
Wd/n2xrnoC5hWvkTiKXbc07pA+st/9/6hoJ1aq5j8lavkEgi9vcHTEmTSHxTA2lfAjhccrCJkyj0
oEFm/cCGWLVPm7GCJTQHPQo3E+QfAnz9UTrQX/q3SS1O7ZLODCsTVqfrtGE92i5bOf9c5JlqxkV+
CRpnlDx4ZLoPX3sSEr6C52R+DaPcLImdtGV2+eMxD0hf3LDps2ZblLgRETzy6p2S6x2mUt9pr5Tg
4yLIQxQzA9Hgal3n8xHhVx27DqXO4qb77DXRTt1Jwm3qoY5NBhleN0t6XK/hXakZgOkgpBakllID
MY5G5WiqHlVYVXIyx0DbDG+gQ+4nb/LU+loti2VLtRylWgXWdPxlg44Wj5C2BsqEmRik1BoU3Slp
3E02Db6cENZda13kgd2ElIwd6khQNGtaVJyeh8mN4zZ6WQq5pbqAUPvCxwoKA3TE77ZxSJ45XAmW
lL1KCgarxa5K6oj9nK+MV6DJQEozho/s4520HyL8VMLcEewkmxyk67z74KAM++I5e6o+yanwZRr6
J/Jq3h5hwi3Z5HFpRK3tgZfOqG/AX7PCSTDcuyHRiGaq33lzfznXidNs1Y1eYtlotXJLjq7s/dBz
iP7n8O5RY8+CWOEHAGGREtRCBATGdOad9R2Z/aQDyTL7aR3ThSJll7Sl+ZdhRxKNxfuO65g6grbi
ce3H4rfla7NUCtPTCoVcDqUE05R4+N3PTPMlMshay0wD/grwqqtKpzGbbW1Yv1/uriVrNSSrsxN4
7P383iBHfXZlOL+bb+tp08V7vTsbZsSE7wrjK5UQJXpCTnPpE4iwMsvfku7Kn3156F5HTdexJzUJ
TxvS9ni0hkhGnoFR9vdY6y0wqcGpGG4Q9gqFcQGrEyj7JEGyzH7nckoprn7+U1YFscZk/hEEj+Lu
2GI/6+H7tzSHCbCo6ZoYN2FZR/hT+oz1LUt7uhx9ciFs/XydyCvO4HAQweqXDV3wsH7pgc2AsW5V
gEBGjECCS+ypx/oP6aunUY3Z2hDgFTyjzlUl/eSVkGEBGwa9or/XeVUj8gCOR2UmzhHoi87AeHO/
4XTGCXWaj1EhOlJE86dAf0aB9tT07cfLK0XutjQTbC2457/vicdE45ONNk1AYm0JKuzzytS3+cy8
5U7+XlZPZDR+A7dTcfg9Y1ZDMGDXxANurM6HqtBCYJ4iTYkNFbt4o0MOlXq/hC1rUwRtW0udY27P
GnSerwk0TYv5xorTXYKFNivJ5sequeo3ajRAukJdq0VwHYC7mjXgh71STNbzWtsdksae1R6KS5M0
l2hTWUK5ae7pjBqFYdnhaGkbEv8/0cTe15LXiNO6r5AOCq9fqhCiAsOGBC+TOFjdQRXpcGf3WhKh
ddTPQc9CTqdulgcH2zYHiUR8PBwLFZ4IjNQCpWzykk+ulyrQygSAF/yq15AKjefmwzQ1ABLDobzQ
weUaibwh+gtdIwwVswQV0usPEzO99uALKWbsVsK/DoNDMVokFFkXhNGwOK8zytxi5bLY8lyuU+lp
mFukPD3O64OrP57sscM9ffgDaBfi1QBXdAd8kLufAdUDmkws3PfLLAGl4FUtAZXC6Zx1OV06DDeu
4cllalIvDfvMs0iWGqbQQiILt7wz+SWg5NFbxQ9UaGoJcvV4xIquCGW1usVcGm9Ix8lZdKHa3jZa
oSEZ+ggasIqpoYtv8Uwv3pft5vJEpGyORDkUXANdCz0GX5va3VkuY7TxGfVJe4ViS04VvSvkbm3D
WZCFs0AopGlusw4JjQaznKenEZdoSpcz0rsmoTzJBKWyVx8je7W4JpMgn+R5W7F9Skz2WXVMFsSL
A5+Afvx/PD1vf/0gqJZTk7MmEwkTAH1fxNDBZthOOJyqUmWfzTovICDmvR9J9jCyjk7gsbbWo7ga
L/EJJeS3Hp8EdvbUHIOy3z1av34BKrnCZK91rSsVE+FjrPXgoge/62VN0aolC3POAqGAoKLo7joY
fz/uIlqV+3TQA2VJK/yZAKSzJ94ABRYtSRBwGRaF5a+g91KiQ5Ks2g7234v1NNfjw5ZtNH5MwBj5
lGpkl+xr0qNQVGfW8wLllkouQ9y8BOCwSSTtkM2d3IeSFTLjIDjoELLK9dMqKmjnrB3/GQmg/1Cn
htPR0sEUCue2X/QnWNqgyXGSsl2MsFJaavKtKhTu6HFmbk1mSP/2KclTmbkixgn8sybKxpDBH+v8
MAe1f+W8fdIZthb1Z2Asnnc7t4YLlOfM4DtKfSrIjYtAQtv+cEjSPUTnu4pffuAdot9hJ8AdOYFs
eNRzlvEmTZ4JWn+cK5D/Khw/LBm4scByo5Bup8F6VgeKnCA/ExyWyxEI7o9ROSw3F6jOFJeLea+7
EXhI8MlDZtrgWV8ktgoaG50jQJjdKJl1YWbX+HFRRhBvCamBQVQEe/beSzbmR0OS5fFqng5Mus3s
e5ugxgJ2EfUOOikrLAopPzpklTXQ8WfDZ/rQ9SD5MxUyr8HoLOZjVNtMX8XiqaGi6TnC9379jWQm
6k7D2LkVHEQSfmMm2JtNwkI+dDo6EPaw5/YTM5dvl+n+bfhlmVtAYPIsvmrkuYUHrPNdmpgMCUOQ
Xo7DZ+2zjAKWAN09jycy5oUr2kZQJwN0hEZtENpA6XE3004z6rDAVuGlT8VKAKy6V9TNhGlhZCPS
9Nre3RiSZ+BIDtBBJQBEAUXSWxwn9Gxk5212ywt3//ggKYZQL01P+dQAFDnqknpDIXE/TRRndPz8
u7WsETUWq9ZcCZU5PXLsRWlL9jqTWqkRsNQQDTbPJDI8qoyqPt/yfqyZzIHmAmDljFdnSA6yNekM
QnGoj5vAOwFUAurMRcIgpqzgQ1qRSjXfsSScRrHEErLzLTLDRfYI+f1fuhYf9WIi6eoi3vVO5z5A
/WB3NxVabjMvnO2w9kxjd/E1BTT0ZA8637hju5jtEDaurPRNhBkjarqPkUCnCDuvcM8HlVVrADhU
32qlajxDml8hhJeQiVkMmMcZ8zxwEAePW9Zc7z9mskMvVHLC3Z+pNH0Dv9FXLGB/mW06gY+vhGcr
9xoUCBylERTfod77ZEE5UA6H53m5zxc0GqW7B8ntB+N02vW1nuBdPb0abBymivlNgZhLuzwPwUh6
SxMgux97Ljc+4c9dRkJOnCHrnvWzwcmsYN7PaiM0d6ovPoVlKGeuixMbcRTyLQX0HfFwIleVjyok
u5V0l4hZsiYXuzC1cup7Xi3ffBoLvc+XbVakFnqHaI+W664HbGqvvzriNKI6zcgUacmidi54XWHh
QaZUv2xYpgfFPoqGoDwJf1CqA/V4tl4Ac9qbwoFHrecgQQGdZUArsFGB9pnVkyVXoUVL9lVqVp6n
ABlvBmbcRp2ywW0cowDABsSITW/GQ7zo/o/arZbjyz9iErx6+BARCEokO0OthpoeJ8byEO4RqNGO
qrN1dhGNbnNOLVZ0X5cWCIx/fUK59b5QDnU9a2sttfmksiRNVQpklFz+ewTbqEFBQpiBXUI33pmW
iVSd7c4c6O8/5/ZvdL2hSfCx9Bb6PCWaPkGLotDikkpxIq8jNjrqzi7K96l8wx5jojmJVA+iBGge
5qTwIAwypdO81+mOqgztj/Fz/W42E/z4lCsP0r/BD5SrO856l2nYZoHgEk5RfJtcHVDVDtdYIfzs
NoHufJ4sRb8Cgdp8l+5hrdxC44NIkbAtdCB8uM/yxOPmR6OSq810UhGiS4Q2Bc28eykgNoEvqPOI
DnFrpgysxmjxToel/jVLztOUQIrkTNqf0p0+OEO31Tz++3GYsSb3pxCp/fJWHQGk3SPQ8YBoxqgh
cDBLI3AGHxDMPNn1TCDq/b3nPaBxKqfKCCzIpwhTcqAv/QgyG8CzaRXGdnE/EKtNvLwc3QRBsFyf
rXgDJxlSYnC1dZabSmLUPYXk8k2ki/UJdxK0qjI5jeURfE4pXUN0X26JLFEWoIPv6A+BgJFhvz0g
+nB/dNoBTkc2rbjHXVVi9eQVqQDLCrpLDSXGz4jWjVnMJ48XUnVhFT+r++W+9Q+e8kqg7vCRULye
MqOe+EVIERNLoJXN8J4qfw66nChJcH8lc9Y9GXmerqSxGuNJH58JF7ewmefLE+v3MQ2FIKcjHAqg
/eF+qtWtiC4HiwkRMww/Ko+bLnWzsuGhIbQnmAsPCE9+Zw3u/7AbLHkekuFSLyCUSAntLSOi3nbl
c3S2kgM7GQHNaGRikijyOWo6kqSskAHqAxbnSz/ODqd2Do+mC+btUviHWZTDylUb05MnnmmJ5Bfd
0003btMCSdWqDxDecVwMENtsjbLb2ujY0pQQ4waQUWvF1gU2slHoaldBjSajVXV1BKd6RXmObGZt
gE7aPo357whe7giZeEe0aQhD7Yb2+7gzy+5A2kKDrzP+MPRwIS4na0sDUIMw4pbgRMTKPURPeTnc
m57QEwxiuR4MuCuuUhSE7qdBgGADEdPF/S96kw8ddlHcaFmWMAgWXVI2KHL/Ypn1v5jth0kUp5/X
rcAHzMlGtEvg1IxU+oG24kiXJ9gCGL5hbHElg5HqRHDZXCDuOq9xD1OOHBFjlnMr5/bd5nMCUfn8
3Zc3QYJwNuPKO/F3lr17S0zNcPqJSjaaD6kXJwyARl20yDIYrJrPP6FMhALx9QYlpx/MeY8uHJqA
lH/Xa76n+XwFyOpInQWVMKfLnCnqLYdF6djom0ynHN+Ecv7k1puX/aZcYYIHnSFJ7ANSptWn75cL
/+JatWqhOK34WEY/xmlZ+CxnL7oZ3zz/hn0Rn5Sq6S+b+lAMU9YxDPefvw5CFJr92N1IiEle+6Ph
2WHXisxySLChHHfXRjwCMR3X0EYDg0SUtdOgYNrEEjYZO37Wq6S23bggq1YehOs6y9rfjWyufLbI
uWcsqXA8rNH9UaaMtEWAwDdS4Oc0khHS3pyk0WJOoSAx6FJhrUt9z/Kqw6uOa1teSFfhgKGK0J2V
+9R7+r5LQkXe988kGcd/mPmPb6J6SWIixvy3+Np3N5AoRs/kcZgJOpBs+wvEirj7kUvsRJ2wjVzi
uwkhJb+X13Zr0HXJWzkOdeXfIB0kvnTdOwb+jr+BrI29ky1Lb+kE5bHzgk2U1Imv8O5s3nFye5eU
czj07F4pMnInvqWNqPBCr31bXgWuBiK8uybJCdFTpl7pSqzxWdwUwFMcGBEMGTe5TYS1hx+s77Gc
oKz9OzjrY7j1eIkHjAzk5JkaZwviyU6MxArfEKc5GUnLYZFNSUQkTFeJEuBY/NwaE92ONHzDklM3
iYpYxXf+dKLdih3sQbZo+FfmsiaPSCX0IS5hKnymTwZA39Lq9GgKNXIYpKkGICdiZ9yCNTquOg0A
bJIbxUSHhTG64CI5EzBWfK6b6KsRU7HiaH6OGXoV9AXsC6GDD65ys4K21/ObaQEqL3W8V9Y0ugUC
Kv/mTs5sTNwSom45tyg65rmZSRq+vBUtq0VLiZj2u8nbsw//XIbEgVAhxFAqFZV6d/vIh1FTiIfM
EudxELJsjRFhKi7kgzoquX++8p9VSxumsNLzUwZh/wv3lHj/K4owCiKRX3NVRmOb2FKL6O2Eabuu
QuOpn9sFSQ7s4/QPXdsLVyoM4MRHmT9LzAvyIHq9L/C4IdDs89kLaFXnz/egA+APpruyvYgnH40G
F/F0Oop+ArT9uNYpwLooou4b+SjeqBF0MdXM0YVF8Sw2D0atsnYmD0cJ8x2rjc99xqM2zVSHwb+Y
eCMdNIW8WT7jA4p9cZjjjWp302ezHGLKPHTt/0KPRF1JaHM9b5hGnMY7Iy/vVwO1FF4oGbsfIdTa
BB47OpgT0tulJ9wLymY6LinJ8U837HaZEcub1zilWmZNJOr3u+7RXBsinYwuuHSXqOUwqplj6gtm
iYil4/uMyPaIv91TFDRmc1YeFFRF1g9HVPI7Ws0QQC3cUOyFOAsazYNQpdON21vnRtgB5SSFcsGZ
QjTyIBrsQtNPojpmspgZmBRoFK1hWaX7OuzzJD4ap9ItYesmgkp4oYcBJCEmR4SmZYaoxhQmvX3N
3aoBrpULVe7ddt31GLbfZ9O61JOBIobiuWE9eawPQS4yfbUR+v83+a3mLyz9yvIHByKcCoSQPcqX
ZlCC0dfG8icwfC5MqPgIiMDyxDwSfFbeEqpqWilP6xefqxcFjt+s9/nRGN6KB/+n+j7SWi3TgtLu
8Bsv4Kg7AIi606aheL1R1Dzi4fGfJNAExT9WWufSbPQmAEy8tvxUG1SU9/MgriXp5O27Qut+sJX4
UYH90fcFLWgz0ELEP5Y4Ulbzf/vQa61uUvA6UoDSxlBXJMeXxzSvFUCZak8+RilGH9o0Pv70SgW1
w3G4ZRWy/xYh403aeW65aXUnv8HOu+Lb58SsXfMbekE8iklzvunLRBjHLu5/ZOoFN6Y/4tL+z0gX
L0w5jsqSLkX0ja4OnFRSu5305OlEkzIaikyHhtohqk5iCt+1+KM8vWdVS31g6fbe1oZyNtMvwy0K
XR5C1HjXRXmrI3R62HpxXVK8PTRC9mHUKfiTKGUU1fb0nUe2a37F14QlacfXr3jaB7MOtanHRgfw
Q88boGw46bIOLzj+is/fCGMHOyA52P/ylDegBPA6zdjaUk/GMG8jENDHOdaQ2Eyy5lSe0Az7yhfF
+liO9w9/6hal3n1Wceh3pWKphE1ovAGAn85WrQgachYUZHNnk8pOBSlCNYYGBl7rVkGAlKoSSV2/
OIby5DfmjmCT0qHxR8WdYfochyZnwoMNiRpTqDfDN4kOcBrVdXtY0l5B62RefSvOjBevFK+rZ/HE
Z0VAwfaFgL+r1aciu0ws1jXN4+Bd9j2MlCFX32GB61IyaiXz5gm0iZHm2VSPYcJSUtrx/iQyqeaw
GTVFVlQsQCLIHUiMa9Mdj/DoDDKzah6PwNpjEgcLZXdhuzXluh52c0WyfLc59/ZtBJazFhTU3wVu
dbADiXKhbFcUat4nM4qD8KLS7H0YoiNei5EqhU9t9Xa05na/0t6wEFCDfTXzG7tmARSUkmI2Nqx1
38O8WbCOCBOyZiO/xlgs9O87Hnzhr8jB02Aol03dr5OynUqjYiab9JzYerqVkoY2UWhCgE1YtDJt
/Og8M//6gOXqBW2YMf0wyT6L1v/ZauGJKP23B+TQJBrdP5LxS52cJ5A5J0Qea3rNoJEqMQK2JJ4D
Pt+dUQE0k/kcFyOz5m07ux/6lBhgMM6ZgayIEIFvTR801thOnz7QL35+G2HjeKrxNDfrnY2xOuUb
V5uf+AJCxKNqS+Ek4JWzkEvwj+EaBaZfSYHjSutXe56fOG0JD7TSGdUsZMpd920QYHRs5VVVEeQs
G0oiaMQKpECPXyM1PQZkj6YkLPiGDDEhN9MgmP7KV9Nrk8s3xUjasmXHAL6XEya/Amln5EkOcA23
gGx5AfviDLqgZqNrjQPKuNZswTug21v0ILCv0lHFqlZBSQTBgdZBsYxqRbmhv7jW27hmAhDNhYM7
CG6qCAEsnXqCJmmCZJ4Pm4OMcl+UAU18SZi3ZxRJdqwqS44mHNuCHJ1/PqEnmTj9wNJxw36D165j
bzAyHH2qvBh4Ke743RBMyESnARUEvsVZJ1Nd3i6Bhfolss6O62JcNgwaWJohIvgpSKeLSxvWABHE
/FrwKUkapLsbSlkfMyzF/xtjYeiIPaonsOCTEzHWMxTmvgaBp/0WnqQJZUP3xYsrJpR6lVWpZkJ9
Xr1+pXdzn1RjIlSkkkngRwSYPuC34mILeHe4vLCkRO3fSpKop3j4ouPM1knsTlmBio7pkQM5Fcm4
4kc17S6CzO24Z5DRJhEcV3c/CKshHOtnVZtTEKFELe0uJcydnq7zaAWRgswd7FlrTyW9yi649o7a
E/XQAqH7uJHef8yAoqjzAPh20vhfPaBBaMDqkoUSGL4Om/ii9RBN99XUq8io9iewEtGXJY5mBsWy
nRpURnF+x0x0yPsR+1Jgaw1+j99sfCh+n2GGinavdH48OKZT0cp+QwG7QhiSYelyE/s8ku6W8hZm
tSdjAdMXQyNFndzM+evffdvQlAJ4IUq4sUPLT3drQCr7V+/5nQ7KjzogzqrYsDb3u+8dXP+y6Z/m
fPzu0hUL0Fn8ay9Gn0JtL/nl9GWEf6hRas3nSaz0k5HL5qQoWBz3RnY11lO07bfwMTgDHKHLQos/
f2msrJ//LXtWaX5OAf+bpbsFypp+VXCpipLFa3iBYvuga0N+49aXIVWsH3vHkJslTUxvqCYODkVk
SHVM0LICHRHP/v6+bGUyxqdjDT59KAIl8t+bAocT1fw+4Uyil39a5m1hcKTdaiuROl/1jgU3ycxe
9fd+xLztO11AlCZSWYEsffmQKCqDzAV0oBLKY7+iAb/WP3Xs4SNynxl0SvTDe1wzpWoDFUuVBCOK
93TeAyYnTf2HGGgs4LXJnSHy4gSR9xhvFbMiszN2hjKjVYuAdgR6fOm9QKM36r9ckm37mPhs4V0E
dWV2vku4jTTf9j5yxhcvEYDGn9B92CkzFnXCSu3hCDVrYbzh3cpjzr9nuFHM9SBU2fWrLcyTWsH4
RVJgfIPz1yIXYc00Irwv+Wj3EUFe0Lf996Ekr9rxZtNdGO7zorOz0gtcAAslib/NWN10wqg6VIt6
FdmCFO2ci9B4QkZbL4owmOwmO492FLMBwEb9OTTyrYehI0IkbVlivD5DeDglDgcfBv2sLaz+/hq2
S/DK3kpD7gRp0P2mCJ6l2SdWQdhKc2dnxwinh63InYXuf/6t6jhLqrbQwOIXR8X2KxB+JEDFEKCk
lt2KwbV+bMdgtNxEgTnyzmbxyXAiRd1RA1pbtN3qq7KawxNq18vZa+48X3sc4Qsx12jwI+lgRfvf
8AFrZKM8slIIVWkzgtgrgRZ8eFjS7tOnoCw+YPLshx6pen6jsli97BLGPc+9BR3J67tGF5Y8C66b
GE4ddfkxg6mKZOBYrerGBmTCnTKR8dw3D2FY+akYLNWhkKHV3QRd4O5rOIEAy8XVRULelF0wvfxA
p3ko3XdH83ScZ45a4y4M91V/dJTHWfXHamhaTww0l9y0zolowQQ6/sByZs/txduQ3+ztl4bXSRLm
uCmAfnqBh47DbSksOnMA9amQbYXIxSF8OJL3ktEuHh3RN7Aci4e6RQlS9IbWnsjpgC6D7yl6ed7w
Pck/mlCf13CqDLhp3WZM2J7zIgiDIOCNXe61sJrdoBogyZcUQNcXl29LZbBzdeRLbTSFI1gqYCRe
U7IBhogxzJOhD4UPzgaoAcJQnGXC6eJjQwXBiV6lT+B2TfL925zsT/vQYS6J/jqVLS+albeCS1Re
WOAdfPxBjvD2ZoCwiizXtC/5FtczEvyv9op5MiX+WtgZkEWxjdIOErrYOSeQyb3rKiUBIKJrl6Qo
ktsXpF/t78ytokgKMVYuKLYoYxWkoMlRKDyQQeK2ge40T6TJseKea17OZK1qlOdeFeYnkpQMeWQ9
gKTrrbTApidSxQQryn7TTh842LHicr64ePG6MPuBI5VsDd2DyDm86v6PYUDz+y2kDyplC+RxpF8A
iIJANn1YKxMJX+SLQqHQuwli6uZxTV6Kw/nTGb++D7tVXCr6pPnCY1tv8tj7MBJNcU/xmAGxqDip
vDDZCA+srUATPL/lLCmaZyVyC7pdMU4HybCOSvvS2PtluQWW8GWh9FWYmVcISefWrX3GwHuwZ3Nr
CnUt2mDp8iHZnC2lcS1ml4u5Kru3sCmdSGNyGavLbMI5ccflBCRhbk4uR8uOsBD336aqDM2s4iTG
m9UeYFNxUe9bgrtOm75pj05kQ7YzHtQsZbT7i0bA5NcVGgY6zRhgHlk8Ibmr1feM4h1xN6xqborU
GWQ03AQUxekTF0YZpKPzDCOz9Q6mpwiZwZwla0EOAN2f1lfyX/4vawwEGMhxSy2yLkI19KOeJO8x
gi0wt7os/o+uYRrEH9R63y7ir/uBRPUyju9q5RHA6+Qj71lKag79pXG4oosaw1IjlhwktHEVHz/M
GnvoS8CLcH3aTM11GuYPUsbcMyQtfr6N3xg9Bzatsmg/vVzIOLajYNnCXJW8quxkq37o5pto9EPT
iZWOyxkLbaTL9J2fAXL0FziE5GsqZqveDvlGk/tK37MAkjAC3KTPWD4EvVFX1D4m9HHCPzGGsaCQ
bT2lBqLdJcRQry/ztYuyb2G1ddHaochVC1zkDkYkaUfFS3Ls8E8UfSqfTYkuatRK4wrfcTM6QCEO
dKwYdoIXG1BZ2mM6XM49lRdNCXjZdLt5MqNmVbPLdG8hi2G1AS1t3j8fWVlHwYpZQkhLOtXqe9uL
JcX23wemfbAvt7stMLuSPO3JBHeXWDe7zyQfVVm1YnpiRq82tnd7QRp8Ludjn3BuzZmXb6mRIWOc
AVQsW13LavLViQqXY14gn7mk5esMyC9uJbfmVSo1MzH86HZcIxH2vNBls5PCmnwG3sUKT0HcsfmH
iu24xHEwqHl3nb0KBfY9GFLqxBarv2/LI6TZ8f8p24GLOoBLQ6/K/P+rI4cODXSkgnAAUO7itt6K
PM1lGEFi2oIhEq5G8NiHskLuem55Ei70Qpupm99ut/4RvRaWfVCWx5MaRMfZk6AOplU5d4DaS69+
WK3r2yjKQtLJtOr7AxeKWP3EzpqvzpMpVKBwkjMhgLSdn4b+AoJ4rUd5j1BeUDGrCyZymosGb8cr
PsuhZ6aw9JGyRH9V2kxikL6bkbaqzpjqTDcMZqfRHP8O5wOzA0BNRi3EJGWMH8f+OHVIm6/b/Zd7
RdA4ABDChuNcBGT2NsQTrkEAjyGjKqxOO7jbUcBIrdBEr4r9tpPc0xovOcoDZRcY+PrDfsEJ4KdW
UNiorxhGtGYPJH3iS/8kexYbf32Wc0aeVOZshmbEHpFGl4WtIc0WgX2V+syTMHDGyn2vefo7dTXq
yx0t6b4Cwzu3gcAuq2IPDhsAeBt9Rwd2sXen7zhn4Ey0acqwRMj36f90vDTaTbm7MryUIEdcTim0
UWaxSuSSXBktKdJmDTfhieUWn09+0zPKSn9+kxuUPVmxpU0z3WkMcyn0TY4O9wpaOkL8QX1Lao8o
nknKtn8rjfnT0pPLLdjzBlQZ6D9jk7LJqKryO1p+XnFG97e3j+y9sc4pn5J2WarWwsaEgI1SaQDe
i5cogQibh/wjWJqk/Kk2tCbtNHyxiTGNwl0aINSzkuRe+60PSapHO2ssYr4HH4Y5RncT1Dy5fix9
lFgFKKtWLJjlbyoCTW6m7/AgGnFLcQpYBYMAQuMSK73rgrbKJyt0HdeguGztUKQtRAegzfKOgnLW
qjorl/uBQbzJH+PTjzU+EpT9voKn8ckKG7KaQG+j0aOXVDpMmdwBdeMYdxBocCSw0H08BsHEhPcA
OzVbGRDkuQQIWOedK+e+83gRlx/0nXzXurNqq1CIdQg2EzgCXv8y9UTzGB8N0L0tof20onqxRsuQ
lCIztfba0XuxJx/Uhz7RtEbJpGmowMGloYwj2Jtdwus2rNZABTYf911V3MbsTvwT1qF085XppbXP
SYaCDg+ycFpgadZwjaOmhDsWMuJX27K+yoI1T/TCWxYqrqnIUfMvX0EbZevvtqnJLSpC3GQgIyvd
zC/eodAz7aBrmj9XiVIr9hdhvRwAs8uIIs1gjhOhcgHlD5kI3P+L66z5W1MyXL/HNZTEzb8j59HR
O+wFdYoAoXfy5zyf1Ea+l1TbgFrY2sqbBP5HyBVLomS6cL8oFs8lbXdSpAhnK1hNz5G4CnoWMmZO
dnA5g6XXvZtMTEmsQfJlTDffLpscpE8oNbHRAWC3sYfSyhaqa24akufNspb56EA9tb7gPMfohosj
sVHNoAiizS68NEBOCN5J5gGFsOVWitMOLrDcgZ8L6tNnx4dq10CUlNth2YtWS/vLX8zydutoqmkK
uN7cZ+q0x4mdXdq23rhj+20elUrx1bCD918clTnEEe5ujvtXnQiXDBn7du0ijnvcgA9c5lEInIWM
qTnlll/xigrH9vlKrTQH4WENZ190kIUl0Pvy/vgBJVQ1v8bqPt32ZClccQwinJhPPUtaHfHq8InP
xXmDf7lGzDnpP1tjTOuaXTLAMKHnMfwstnHdD/V+jNgAeE9gC+mgrctEbNtlPpktc/FEBrnKpfOm
nB/fVMN4gRNBLp9L2Wanku3ea51hl8DJxCVLHTBTklrldIbZDjccmz6E6Ye5fFiJ7ZqKYPXg1GHT
sTMDhgCWNiTcScBLzBz+/N2SXgNceUGtB/aW61I/2o8u5rB7ct4IJQFd+y68h/3cTPWq7GiIsuWi
fiGk5zdqknGOi4XGZtOPqRZkACr3nm6lKw8izvqFUQy6Ei/9nDxKgeZedkRL5VysH9kVV4W6vs1R
RUZ8qFd3UZyPLUQpWsIH/MS2IOhBufPaHfGoAu6x8rY0w7wOXlDCcIyK0sPvl7H6KGC3fVEajIsU
8LPn8etarCfd5rwQ86k7svbrxEo4cq63iabzqPV+Msb5ohEZH7cBdWPMBfvLzwmrKtFdWcA4wNw8
+iSZrhRVUOnvV2zTHhvcpXZEZwJHn38Hy62AHZzFC5aBb+xiBCnuYRhFupzl40OFxXCJ9ay33o75
xrqcpqL4lRGGniT5kKkzkTh4P0riFlq2RStsIpoYHk1iQSB1IQOXALgJBLMubWoG3ZwCHucZF4FL
CRfKCZ/03giCF0BgMSpqYrfCI0cr+RmPWjxnoEZVo+u5oZ+Ra445Pdx0KPiMg8vBG2HvKDpV4/5l
kc2nOg3PhFBROOanjhHdgslHYvI3CheyFbtII/HDVWkHZopkl239BSW1sNsofP+vKYinUO/+du7q
JVK8sbXtpapHyWf0byA0zi6qGRQcaeewVqkGPtQJXqrOIgGwRHY1EpNIt6SSd//yb2q+DluuUeCk
5+2mCX1DOHDfvxIG2PJJSsjiZIEnu6442ZD/+yxeQ9GBY+MtotIRIgPWoM+9RO3Ofe50fpju1Ds1
W5OH67Xx4pnONnyVJK5hddR/WUOEczFB6btCBWYE0EJAI0U9/qEZJAN4SDO1OTfPMAMYTJ/QQnVr
442PEow36m1e+SwD8yWNKVYbLSoAQkJCSyGvDK0oraqpMG7DjN6E6+GmdY6PSqA1Lhgo/bXyVfEr
96vHPjp4h2Ksd5j/840RAGSR1G15YOdH5ZkXj/m5XoNrPzCHUSV7wyh22KyRaYyCaFzj11z2y6n+
HwRGf9gjcNFweiWu2keKPn/2Y3XuVdipU0IfhwSBtaYjda4dHuqRNx0O+frEpRDijJ8/v1o5wAzs
X0gx25hCNXyRgBBKj3nQr/5GajJHjvIBUmxTD1sBdVUKXyVfk+WIu9IUJoMOk2WE7WrIc9ZnDenx
BFDkxnpXy4OdOJkWpjzCWbWN/yTWoMWl8Y8Qfck2TCCG5m7/QvEp26KpApZiWoNWwJOT8rugO7Lh
PAgeK07uvhgddI56uh3VUcBOSHrgbqFA9T71V65FytfCg2mJHNYBfJEFE/zUKE+2aHvi4gKXUHSA
v6wq1tEwml0XLwZhEcBJOIr+c/JWMP9ul5CsBoDgyBbePQC6CsXsFy3WySNsU6ePoy0wecna7OrI
GBR2RTk2F3C+TxpvhtfGEsV9PGMF4uQ9G+I31SN9pRqk3Nl329yoan5AKMNP9BCHuzSeOBc5SZot
IvKCsO/ytGj0sbn2B/hu5gwKBG3EdjkNJt0kodeL2ef8+aewlnelWV0p0xG+PeojVvOpiobVRMCH
Us/ZKTXSvmP4KPtGd+hIkyESYkFf47Rqs53fTvZT/ZnbdyFe+I0UqXcghVsE4H7xsdmhDOc09uWJ
EU1t7lFe0kDn2+nXF7KfaFc4GxX8UDSxDDmqQlBrzrYczwNZpXaM2pUPkb5KJ/00lKD7kg6WqFRS
oEbbD9ZX58ZE7s3Nud4cqPkhVbvz9K+ZDaofvOnoDQg5USa6WhzOFehKEjYESW59Kfz4u58VY07V
RTQl4wJuMZuresYsGbARmXkYIoJ5SGDFJfcVCIdqkwFlxZPWhE1ttxkrlnNmO6i/cvHoJPuGMDun
fouHJ1TXouhzuRt4eGDXmIC6wKimVyaadPbAzu2v7NNTBX7ipb/SNKNV+zireStk8IvTPoVm4aPJ
HglkburdgCR52Q60L+nbQY3PZuy4NCWpV2pYoltPuQAqD7x3E98f/4o4c5AzTij3+Brcty3ut/hP
818x2Xkn3pP9XEWG8Xsm1KbfJbN2H7p5NOKwp4QAAo+lAlpdOUFlOc/fHwn/ezXlxytdM2GvdBOM
+gX4TdtZqZHhlZpigyy49vGpe6UVW+XPkD44LIEtKld9bzzwxWqajaOE7SvZwWs3p6HOAZ+cqpCI
COLW4MME0FI8IdF5dfdgsKnmI1boOhtbowFSRnNWXbQ0HjtrlhwQv2U8rAXiChBGxNv5zkwlk3N0
3nEbrnt8xFgwp3Vbr5B6u/siwI8KimZfU2GzQcwvAw29eKG+gKf+gGstgpMQsr5CM9ehlbGbztQp
ae1kiXZopuLuo+BT+hAA1nndV3Oo8t2Axanpqg7HN78MtEfYneSuwIBVbzTgA/TLO36awHjCoz5o
Ik2K125wudP5RSt4+2mdMreiKnzDF04gcmzdU25eyVl5H5jDHf87UZ0L8mSQBO8sgHDJJg5ueGIf
ZOh8MlnUTmGkHqngMYL5r+ZI2J+a9W6hJ6O+gKDASnZ2KOKRCzS7zlZRs0qzf6pLGuJmO42EjOXW
fq5sZHO5r1dDGkX72mUZdS35jD104dX9wYfKXt4yp42WiAEt8MlGRTAYmNl3rmFmAyHErKOzgu1s
FyL6hWFilSDRh2u4OG9gVzG5mfIzVFuS7acB5ofV1mkdECb3iKmivIIcySLQB/rPbGMuggS3zYOB
Of8vyU3zsJqtG6a+B5f5Ur3X0ITFQJAWpB7IrbdQvkpjLKzfo8v4bFZ4Aj2znarttNieaxXkbyMH
xtdl3S/7UP8UQ8xAK1VV58VfOITViTrKTv4lau529StC5z6G+ByIaTZpA67VxcHGrGIrP46LpEem
Lswv3o8Q3JA+E9LTCUttZG06mJ8ZZUQWre58IBIJjtykyCcvjTmJYfQQuoc6f4qiG9BwNyj+iwJH
rZxBXuwgjJ/6TxmIOgTRrzW13KAy3JEkEuN2ez7PUbqpTu3JyThHRy70UtOmuVxES8Ivihs3khIq
kvN9hdeScEb3JEd/IBYwF6PxvZj4odAvGQiJXODcuJlhq7kObQnm9OAdqQPMBBwUWZNg1qDMnx2H
VlXP7bYLtj33RrFERknyGS0oUh6DiqTEMkvnoiwmbRe8bZWdMVr8MNsKZK8KjtrApFQTGiBruAbu
VYGSr2HfN49HH53nM5PPObgn5bPDn9dX/1hEmkcFACN1Qk7xsnWW14HSIWT+AjPT3+NpaVtJ1C85
WQ2WT5igO8Tnw6X9U0w8js6QSkZmIdqQ4O1dzzD25bKmTuhEvnOA6Q5Fi65dLTBxMYtp0PLIYZGb
QAAMFEG1v2Ti9yqMTw9MD6n8TdnPqm9583B2m4b3hkl4ANRhqLch8xVV0oGImGmduar63dpqf9wv
OxbsAkbBcjvBklWEC+pxHCKL5K5yF0JA/I/dWpTZ7rKzpz7hQVYHXCwKp1kbyfOPmHOrunnUMevR
tyEY/PgxuomZqZW1//hf891R1SXaUyPYIBBtyMYOKUPouatJgPllyFvsUb+MV8Fdtr6eOSE5A+kR
zyfQwYbXgPRvux5eJo57uZ5D916iWAL02ICiEz25feMksxrVD+jE4cTIk6DiwO8tFhFHW8TIUPj+
I+4XvP6EjnODLv1iMimgAnUzM5WjpxwPWc0QIpsO0KPiFkqFke5NtDtgGrUo5Ecbwcf/m8jEqbmq
hDaRkJrlm/9+7G0l6TJcydCTIocmBcjSMLfc8WQPuA3OcI609Hr+TWCSlyVH+JguoovAp5oWmhuI
7lVz8u7yVCnxECe2M8aZ7ApMtZxhjBmQGfhzangGxIbr+IFxEg91hMQhM4OlIBS2rQUjIbvpYxmG
Pep/qN18isySDijFxwyf1X9ExDq32m791J2mNni9evBgw1iBbqxSFS3Rgf8yVKHJDMB/I0UtEpxF
sZISAnOcEdnrXLMEQNsRAgCTOgAe8RAFrsge1U2Q0qxx2zSQQ9BT5kqz3cHr9mBg71l7BZMDmfut
Xy1cSlht6804u2shQOeKa1bJjG2ilwqGwZs/38jGg5MQK2FzeXcmNU9kScYy2yf8zLHq+/XXL4d0
jEbW1j2DCS4H66aWtrh0jGSWnlD45B1qL8ILuWYaXPLgDZQBBzXZhhUp/XfKHLas7X0V6Qc+zSVe
y3BIRA/qsGfeFSGwmTLcao6yE4wtkCmxGOkIeRJoXZwCxx5vgatfiu6B1a8btiXRlg0X58UB6ola
nH9YMOhZHGLHFJgNydBPsQ5HPsrdxt+IdMr8pctzuxm7n22duacPtpK9avdvTEWyd/OqhZjQHelr
1pPRLbwbvqcFvCo5bCfvEvxvtLfzZq9ct5oLP0E7u7wdviEvEMZTz+fVzxi/b1xjK5UqdOKYQHaY
KYw5kxs0Xj6ESZzGsCx8a8f+JTDbNB5txON2zB0XC/iaJj79B3VH08JG0N8e4pxjwVa+9Ml5hPEj
1EZs4ij5K8dvlIhxaN6+BzHMEKP0hnlUJFtHz05yVkNFSNzIfxHR5NGQ0a2KbyhINKLk39ab0Rt7
6vRwpVP/Ni/v3susxWhIShH0U/VqmK8onozpiAKownNr9qROOG8GCy+e8Mb2KXRwRsTat+8qC/DT
QhnTYKnBJkx79Q09CPE0iBujReC54QfdK0iZRkVvisLU49HHD84OjFNYc0ZgFUweejC+LyGFMCrp
+56YgzsNaULR89qsHs6lfnH4wW+6QslS1BeHlti7DRzf5kZWuIG4ulBIEw3bhqh8kE43xXbZjva0
tfDUdsFxol2RGKCUqfN8MM9C/cagFmhg1DUyLVriHujH7+N+pG2WUZbf7a2+Ku7a12BwOams4pHZ
4VNq8j56yP5yEt+Dk53eI6jpjqPc8mBlaIngXPYGD+8DLBF3HcQPPzZPU0i0OPjUG8e5D6BT3Q/S
veGT/QvGisyh4NX1PlhDKnUYG5NZHydAE6+nwr6LLhJL92n9v6D031x4ixd1QJdr2ROA+z6gaz4c
hrqPD+TvPDpDgKvdd8ibt0u8oONVU/F8UL+KZVph32EJv5JcEMtc+9ap7X/vJ1N+A9HQ7nkspftQ
CXFt8vFJzD96o1sPfTfkRJ/S9Q2fj9Byv+xxYp1S0FELPhhUFZ9Zj5N4iIrFmZvVSLVfZERus6LB
534OThojEbBDglyVtOlag9+mcPI/JeEoN5HUEI7UUR4Uv2AF5LrtYt+I7IoLdeuT0IIi1x9f5ckX
b46m5TI6r30pQgn5ODc+bqxLCvA8204uEO3o5MVQkJ/p9EtEkMMmsNEmvW5rSEh9XmmGj02J/G0a
XhixtrQ+PqX49mNCM2AIP6LJ/cMYFEJbT+V+s/cjsHyHECseuXWqFl2jRZX8uswGa/9bhoAFuLgq
5d8/R1duM6NiLG5aUKZxCm+lk4ApGR52J4c4a09ofhC9zmg5euzXJRbZRKuhucrNRuDkKLUlB/VF
PorzVI6nAGT0MjprBkCYiLAaUf2aFEN35A6qYDDu27SgJ0ElIL4AvmJcy7yqNrORddgdfhp/EL9T
9cS4pm/chZgsknfbXlC9Q5MAC7caGnH7ASLh3rhj+GljM5xm9nYUacfvK5pqqHdkOXX7r1SQuT17
8bomxb1rOAQa8H+f9wKsn8FvtUejIGwnQWACFpX9Oc/HovlAsFfb0fmwAAglvLQ7ZfCWqsbnNfd5
AWfKGkRROY3OJzk4cLgNI9oNlZb9S+zez49wcI0XEXHz+idXFcXF0Gd7zbp2ANdMfR4nBKuqey7d
aP4vvcbtr7KCYq0ZPtTjZCPEcTybVh8m/74YxHdiUKs/SG32AnkX6g+apZsFETJfKs91mTQZeAF0
gazPnUe5awJi4D/wRYY79Ik1ncn7MmOHLNmOQie4U7vFvGQta/eLR3WlwhtrZBiuISi34m/js1r1
B4ts3QKdzFXCaiMKYUzV8hGfu6W1WwQ7gXx5eynoQJxGkjT9N/wLS4lVm975MLV9EnPj/bYtWxPF
INOlB52eP1TTFTNrquQ+NjH/a6ZASM90dPew0sp+AWY/z3aFN1HCzY9ozlPqh2McMucK5Fe3yl9o
7M6jXSvSJd/PcEWYA+O8cIuX5lDvkRoOfoggT0Zlo5/cEaZyBFGNkj2k11d+eNmwmNRWjk/c11Qr
EusmB/IgfxbhyScZr9wQbrij3OjRgayQDeTJgrVGpbo0ikGxJKVs4jzXIs+UZNoSOP7CLpG+Hz9J
xWGmbUgHTAyjKczqfuICr5ZubDql0PmRqMhoWrYs8J3adqTHIZJBF9Pue50zmQ7lMI15HVe5sL/7
O8MNP9nUH2rmAILNbp1pTDA5asc0QufrscyTZkl+qktNzuac9/FBXn1N6oHanjzRZn49XA1eg1Rk
1++bfAyA/BDvckruSGl9tLAsqQuf0oldGKI5nAlIVnXew+YeehBUKE8zni12Jy+xqJfOLTihg4+H
8+KQ8r3y9Vle4MycEyQFg+Rd7/5mcPkiCzuN0L+J2pJAUk+v7o7ptJ9s1Y6z0pOR9j82r6N/Lq6V
BlPApDwTRh8SaYuQt3mlg2TB0GZYR9UKipPACn6FRc/97vacxXHrKuNq4CdQcVMhCqAVvKpv4IBp
borIn0iPn/hWFkHFBIwZohgNc7DhOdFmciJOI5FljLT+CbFW2cnknw8Ia+zUHM2F4Oq2WcaJM2CB
BcANMIae2DZYnSsIwNCo9QDJP77JouwA236bHgfXzCIw/OcSPOIftkUMi0WnpGvQEq8DOSbjPuKT
obBve7lP7gnk1luHah4DCZS6p43T9XYHucRorYyMguD0ao8j8Cf8zewV5A2j6998ViP3p6jxkBIY
M7apb/9PG7S7QuciGI3+xTRFhjy0kawISctP4wML+LNayubdUHEZ7tPIESEdCXuEj9Kobqq5oIko
PN4Ds6g1vqVy6I1BPK2KawiBh3rD6rVWtLTTPcDQLWbGHFSL/n2VlS4+MlQ5KJAFFSOt/UD4/SZ+
BYRyAmP+d+KiKcWqA7nwNh4V4dplmHxQsdxiT0oSZjnrYXM47Z9whx1mTjs1qe9k9vPCkk3BnQvJ
Zm4MfUgJwMEJ4MWaPcPZkKqoUVmojOyWFBdXoLdjVxonBjM0E4eBawPLNzsxO1LVZdmb/FOZA0aA
UZoCuieX4gwff8CAItGl6QHoGlREcCRjYaru6ly+ZWr4DDUf4DMrgexNHiCyk5c0fTUurwKnAnVn
9coS/7wf6YnlRfX5kfMTuD0QEo1J+STpBT7TBYTGx/xpOsPyWfX/Vv2MqYf+Ti6Qlp1WAauFoYoa
CBUhXHxsJiui5/8v5tm6uXoRvQRv4a/P9YzDpbdi2xxC9C4N0gVocoFyjf+6XyxmqzjdRXw6X/zY
be0i7DRGYpKDK0W6ERvgc94L3yn75kWBik6tw5EBCaL0Xt+pZMsGiKsJxbertvQul65gQtSOnSE8
eJchKffbsNLwcXhodkWW8hOIewFYCB0pM7ZjfaVCjpR2gyiNEMzj3bI9MI2AXZvvBnZ8zvj9uFZj
FlU5a1NUIX52thso9SUCN+09OuVmDJZLVeMfi2ZBgQorhe5kpiGmclY3fIxPfVqfYlb/Dr80LIAy
U271HoVm88O+jaFk8u2jayJy/oelHhQre4eLBpPiUiQ3iWYKecejxIUhbERLT1CEyaOFnhjLWQBh
KY8x6+G6ss96B5TaGenlwsSEmMYpHFpfo4ojky8nwhqAmkHlDML1Z89RM8l1vD3N4vtFgGItRkLb
IIFblEDRUMGy5CU47c1d7qCvohYIjOJzUHMQvd2lKLuKi8IUQQVbdbliqykdBFv1dq+5l120cieI
2/GqL3NACviUhBsymxOUJ8xNtW1CX0shWngzD5AjOIMytwT7K6k53UKiz/vieJjovya4wNRrNt4v
4i4MouoNdtEPHZBU3UWYcJQCN2V0SPGTEj+1H9XT91mQPRyxhkK/mBSw8QHPePqYJVSHRzDzXW6W
/08D4kxK1KUPNotb2TxXmz2pVDXAhdkiYqMOG4s+7ZCDaqdgMAt7xObVDycDIGA+Y7I7aSEXuomd
5m7ZQgikC+RYSbCOmarOzk+tJCM7jX4fYQ+pFp92QaQqwwYHyyPDdhWCOZ0NMLoMvI2KwiPUpW7F
zv+MlHw5vj/DEP3cRuLgIo2GHIfAm9/g6d+znZFVUuSv3lnWpLLBBcjRsiSS5jVS9QKj5FtaKTzm
iOy89hreBwilP6VvkIjZ0Sg4YRESOe/0/On/vjB3WaYXDmCceKDIIlkkWGY55LlS4MA3izWBPNfd
Tb1XQT0K9qiRUErU7AfLscjaD/YS/yG1EmDaYEb7KirPGIFPKZUi6oaUXb2YogTJ4WTrNG1LmG6M
q6G0VBle0tKyphGx8FGgguOZmHSqgGzKCIhP4lCkqXMiZcQ56r2KJfIK7ZJSjELmrXr1JqhcTZlH
y3y/Hs5FrftI7MThjc9HUPfky8YD0LCd6itkMfHz7ElnCswOOWdfC01AWCGdFGNp7MNa/MZfK/zZ
S8gX4xIrUHGPLVyELeoq8uQlgiqEK8S6nDuHqX05RdBr/1rIsrVO8eMv81XYP3kgnUYekDssJ2/E
xd55NkvL5EDqeosTVPstwC1hFnl27Q111UuFioRtMkZyklML4bfmriwMmdBsK4V6arOGyyi1AW3t
fMM2tfGSKLT5HJLb4u7Yg2t4FyzidEK/65viNPeU4+Kbz3ZuU1jVqnDQ2qOBolW0nyHRLaQRzK5B
LaRB52RUg3ifmwUqCo2N3OSjjSLXjMxCQVdF2QW8VupFwp4bNbTKForDryOdv4aC2hb8rgT4Q0HL
YQDrtBBfKjpNE9U2F9UQ0TnB8WXYYMuwqZq0UnHYAobXTTmDjnCaIOrr5ArG91wjePiTNwNMFd4S
UCBshpEDt8Rs9G77EtstjTJ34JbKmacMw/FUZDii6LjUW2AUR4vlK64G/yUgU02D+OnTRJkrhsKd
iuDhoMq0p4SiLXQpcl5Xt5oaAL1ao3ci6fUw3JcfBOd2GV0afhg2ygZfOahhc4C2F11FeW+O41PG
Ze7r9/B67BmLwBB6XXeIiwfzPljajTqf8tzn96a5yxu+S07CTSaBc8x+zR2NUyRKDigZio4nkdga
cr+jBhyiA89P3LhvWWLahuxQO4CdneRB+OUG0gX2EZtdz1ZlSsStv/jT6pjw75ANY799MyWa3Hox
UaCURBy1qyKOxjrW5OX677O3fYC9kIjeMtJq2bH2peqPok/OL3Bkik1FM8Qvps9qrtVfcqCoEauO
zSwUuUb9x4qm4HnsrsMnf1wZvTzC3s0dp2wDB9ejjTcv8crp0lkySdctnMHA6rG2OXXd0F69fM9q
esrJI5LODMcNII5g2bqGg2zME2pEGNVXNFh5V7SG0tezqSVMMDwsYj67yiG9YEzowkZMST++Q2PB
BjhvU6m2aNEkKmr2RC465SW1WVeHU/I/sQ7tUT11jU73lgWDwBPTYLHvM/KfpoJREq7SV+JuLczh
BmlsXJNwJqZH+rhk3+Dn4dJPVv6m3bYvLTB3z8ClgLuLPTsdZe7MGMXTJMyy3jBLUFU37KsVMEl0
IrqPj9ky1OzaVlDaaq4UyBjwfv+SNS50iojhLPeWN0ShGNeoHmzfLGg3mgen3elUMWo0zC2tE2Ls
Nsq9ZDHWCh9zaV8QZOQJDxL/z++h+WM7ZuwrGHpFX0wdaqoni6Yat5lQfoBjrsnrn0QT6sb0xn2v
qd5Ygvhnze8OFLiT//2cgI0JWWdVHuBMKaSYtigVq5j7sW+upoIknlDNlv52KncYnb0ueqxie0oA
u+H+R+PwgRLu2bzjewSp/JKQpbnDD6kNfvVMJp/WZClPnJzTLINCp9ZXX0XomNhblsVIwU5mBjoC
Uxu57H9NLcI/k8xbA2G1mFMPYtfic2ktQtMbAhLgN1Vv53rvwdDZ0FYZjFtFZSmUeSoC5p4KktpQ
qI+Ev7rnP2kr5aKYU+rkfVfOKb2d2eQ2KIktFg3nHHJRt0Tq7GrmtS/0CirbOsU/4EX2aUerQ8um
mnjJPfDMsgeKXNCRb9ssMj2lfeXpHtQJQ7rndaDOyZkRHwjPyBaqh4xtXPsK8dhk86m4Bqw12aOG
wKqWWKK2fTmseNLLrDw54d9WzmzrnkZNvuwSBS+DbQA+R8TMoSGUe2xMCUiOTkhvqNdWn6uWhzqA
bnhl3L21fK0sP0/8pg2Q0exNgkrgaHmvqMTegWcPAiboQ5iTjP4gq9UlbPIaM0/NgkFv7Sf9QG/a
s0wasZ2DKIOsoYtXB3ysxkU17FGq3WPXYCi+6Edu26zIzgGJ+XgIs09RBJ6cyK2R2HPH7ja8laem
zOgQ3eBzL0cmi56pLen1SwAf9ilX272Y7bfpKmCnkPHG7SZnHHaqPOgKixZH6wF/QpOJPi8p8Ceq
abmS8/pjOECAb7LEK1Zq5W/pMgDXT7f8g8fKYnOWnqWbrydvIKpbTmwWfBeUVk1SxqOQc9jubyvM
UgLHPthLeSqzFBdnpNvOmBWdossS6WaW6LNy8Xf4TooTvVhWr5P+wS7nmy6Q51dP6bCbZv/o1Sah
jmfzcF0NVmzKa+92f7faalr/5yh0x/iUgrzd4IpGhgINgIu5k3EOJc2+o7OIabZC5lvUKI3TRdF4
HebfWraJD3XGdLxwcrCG/amPk67VN1QlWE2o8U1GmKTrU93wOvxUz19YxBAZJ+FiXtU63DUHca8f
NuyycO31Hzlw5oZMlYg+GitGL6/PJtHPWoLeGznJP7LOJuC2Cacjl97utcztwUeKtm2PKyphGFc3
MJ8DR1HU6aBDbrKMNxYhMCwGot84Z1NTN+tT1Pmf5tllsk9xD9fuCE9CPikxGwNjKckG2iAFnr00
u3cWaMN+Jye/mTRwMjPBJ/vsAwI+ZyIRdYts9ulFGj9AGBAHtE/svZTCbElF32de4hci65ej7QHo
rgN/DdYrvA9OimG5NWVAdA3PbHKO6OMbepioqlutfVnTWZXrAJgMm8fl5+DbWrTJbECivc5A4FnL
lBTx/eEwoWpuIdGGBqzajTTS5HBj9JB1mMgmAonJbNG8UJ23rJ2R7J/D6hrcsrCRIlPmU5ZzvtBr
I5WfaOKacCBniLpKLUnKxfwl+IGqV/Dc3cT25tME7gwTif9ae7PXHKfn/Gyegzw0c9nNbWFezvBB
8Bp8kloNIGyWxErsd14OdoQMGWnaKJtmZYlDIyUe6oDv7a0Y8ZY41QNE8Pg+cjIKxqRJQFCwROlg
A/Sm+n2xLIYVgDiS6YVFPZQhXE2KrxNYjKv/2QAGO4kdJmGQxZMUFEw/NnLA4heVWY9tNhf35cEH
55XEOOzpr9aq6lQjnLZbLgnruPGWoJI7/pU4tXthhHd0YUWXCM+pB1gbX9q96FeGbagkHpSNcvQ9
eo3Z9VsxSP/ajbU0YuAJdva2KPbEIDRt4dEThFixKHyUcSlpqX0Doa1XxnzFrh7Tzkw80pnhg5ks
A2GMuAq5wNFePtZIHHjtQtMSokNXCafDpxvaHqXXobYDa999T++fuLkClQzKHHT2/yhkNc7HYgJE
hdjoI0gxL5ZP18fi7PYn/bg71OtHjmJSRKLqng3zpiEOXQ95hMJrXWzw2M83XQhNHRRVzsbrXc98
CR8Oge/DWCGfKSvoSySe/+Yr2+y0IIqZXEXL5PrZoCnbA3LTDiTOyaGB3evrYenO3iJU5QOqiUdR
VAT85p1BQs/KcAOX/1US4fuhpUca6S1umO9CQ8sRoH7Dm9PRTH1G6PyBWyQhGyAGgdX0u76XK8Qp
qZNEOi/4hYCxJsh+eATbfTHGULRpdMsLN9Ts4mkOhGmZoF0wWIjclrkRPQr29rJfyLrp6VDzeCVa
9bFl6uVjH4DN1c1gsc5Ndd8KGTifrD8ij4kEeObNRPIj8f04iok7nmZ+CNYLp4s1caflVK4OHT41
LFu2jKu68ekqQ4YBeRoZwDXRLM0lYyQTNt97zUvEW45DjkBeydD4jubkRHNpW8d2Yd503MEkBrpD
K4EQlpTq+AI8TS241pQHj0NVR3LagOHvSviWojb3hSiFgR5x6XzqT3KOcfqOKbLCjxyhV0LEaJuh
KCxrkQFNGrtwAmtCFtNpYklro/vZd+rdjgvOyIIqlQ/UWM1jWoACpTFDnQDrOcQMEgQMAImcBccS
amod8aGQnQV97J6+1Cw4idisGxnctpkQX3w02pyxg0S24YD/0UDZUm+i8vW1ZvSSq50lMXtUwdBi
Se5O4j5rwYMULGvOC4BdKKhINHNjo5JHnVQ4/BoHY1dDD1d07g7p2SJPuExeyMiSJiPSOaJ5xucQ
XypcVSq+UiBMlVERgSHy7Sc4XD93bwgjN35HXzhEzL8htrjLuoffgzz1OzgeTGR0bypRTEK956BD
wKHWfxgnzP7kXzDnmC842e7a5mr4g6FZ9E4w/F50P5CZbwbH0BiPBRTRvDrRK+DDZwv6TuZwWVmj
R0+qPZ1z61vxUCM7snq1rBYKlO6Zoui/mtv0Sp5GG7+hxPm7OnWdiaWReSjQQPjKv3foLiz0+Hei
LohSCvQCe2xzDdd5wZo+R7phPfcXy95G2r7X/fcGGWI8yWbmV5IPjEqAiO5dAEY3/jJjZzHoBwDN
/7lRhXV6OYjqdafjNVDxxroBrz3nHFucg2d82LYoLshhG/PPTtoXSwm41yO/8+8/B5ALw+Q+pEMf
deuUW1sdHDWzj+voIaqSe2tXJiH9t1y6v41b47R0RTdhsoweF5Ik6eWGEFXAYnrWG5Z13sZ+5BUb
n1iA3KWfWgdoXE94pySa/pDxC4gH52nb5CSqhu35Dv3s32nB3N5Hw4+W7mnhm+vkqLAg6B1oDURB
U69PXba8G8uLUyy7xmIOMHBSah2cwA21JDdU+xcTYO67/2BYdxNKZIwNeXCeFU0EFFlQe8h8e70m
keVf4+xFb7yU3rWWYrsKrzgs7EmPSUmCFPEaXPg3jGgrbKa7Xn4ThdO16krNPnQZa9Dz7hZMb96i
UD6XIjHK6deMatd2aMrwb1EnjKEfvFYEcM3rSdXKtSysjmgniO/sabPth6g/ZNitOosNmmiYmXJ1
gmKG2/jZHDB0TWjVOCtXmJP0xPary4lpjse5xXM6EJ6u1uSFT7B3RL5+eoFhwbHPlhguhGdTnk6Y
G8uji5hHx1LkOFTjgTL/+VshWEJkOu7f/jUxvtw87j4wvrpMuVmRLZumjXOIlIrEQK/oMv5sTXVb
glyErNr9Vh4W6ULz+crSZpO1IYRWvLcq9KVQZ5FVSBgJAyerQfeHbEo3HcUsE93Rf0GmVKP0zJON
wo8lWtuROW2gFKYR3gtvTiIfYCyAOpWJyrEj3CBbZJQZCreNWd2H3PCb4gYF8iQflxSfRqVzyfBb
MpCEBAkHXFvXvy54GdFXK9CV2r7NhNcd4PhsjHy1PS8QfArc9YSwmflgB03Ws+idqdiiVDaHi99X
PolVax8Ee9jGjGgkGWi6QBkVG9NXw8S7tXdfMp0970q5rtE96xNlDSu/7jUPjUL3zOO+6O024ziT
kdXNcopevPhrC26c4SrWFa7D/GqqYyJYrNS9PzpbFrWX2eIFJaEvbs+6HlLU7ZIun2tKsqFdkdxw
kV/+jtHLJ7zNYa2Od/tqnPwmons9y1nZ+MPImuTi3NdhVOKLU3dow5I928iXDoXCj5cV1NJZ/UWy
E+SCbXdoUtTNhvh5SwMlaT2nv6A3GilToAridxGZy5uVEm1MCYLQmXSXxzKs/3UEbjJOhrGRE+/t
VjYdZxMdgyVtHXgRk1a9HdG8K1/oa5U4P3pz4BN8WVEPLwA7wi+gjpCNZKEMrgSS91XeA1DR/XB5
LBW7o4SeW4NDI4HNwMntV4YV6nBqFDKQ82+mdk4tTqM+SWEKkgT2+pASb/Jd3IuPvm0oU294dnDe
Op2s/dXthOrIPCghWYMbJM7ZGxXhl9MonyKl3G1fgst5WF+SVGyYsLWKRZpWoh3qFVJtEAJRjY1B
13PtHr2mml7IcnucFcyCasWW9oCsjWqssoPYBLbYSVXMAjBG4/bRTM6OLvRnXqpsJq2ou3gpuXGj
TiicYbFsay3HbweqCzOWkX6FvKd7+Sg2nftpSEU5gnwprfYR1GMR1V0u6MPu1sQM+owUrCmCj8Oz
ZSOKIiuIy4AHLIdp+hqTGRPAHJWwGZP1I9HH12YKiUhr6Q5adM8LxXFOMeGxBCVrtm7pHQ4BJ9Lu
Dacf/ZU6ss7OFFkzbi+xlaSWUJ5lEc21akzwy+jObRmymvWvwVVG/1tDlUvVK8fXwLNnypEsWA5u
bnOj+zTdUYYWP2T9Ezv1OlLZ0gamm3+gG3F8d60o/MUR+blgSQJgA1ym8Gw+c9AVVlYT0f6Z3vIe
IGLuszX4yDJYQ2Xh0zfqOz2ZSJ7Tide83i1RBMLav/xw00MfRmpgH3NGnPSCutxEuc3+GmO/4Djc
KrjBnFye+uMpmUCzqmMPQ+bc4DKN9EY9Arybye33R2LDAJTeQVDY2pErHhEClQnVeFueJZSCPyhL
/5BfKe2tuJ5aCNjXEvl4/cWQlryenIcwkte1QfkFSe2hCITBG7FcaoZ+rG6hqMxZh55L8NIvSTja
Aav4o0Ex4bwvClxk4hd0XEbjuqONVs6sf5IsKhT18rrr+3dcNjQPezbO2BuQUT7KIce+Fs+7v1SE
yYVlYSo5hMN9X+en/gQEsu3nnuS/TD9iqD+2Ir66KIaLRd5jmA/yI7rc+nIDetRiSxcru3OuCl+j
DQp2HVsJOlr9Ypr75J9NgNuyCLuN5r/j8L//AgyzeLNBS9P8g95xqSmlI+oOkO8RO7uUB8E8G/5J
on9gA2bb9N5c37YXxp/mg9Y+79tAGzgG0oRCr9pFrJVgXfwbzJsqYjXJC5KBy7Ov8NSkysVAi7MT
8/3c/OTr2xZIfmI1Qj4fzkTXEV+Y4hOm2sqKPIFrvlBJIZ0jHVDcbLV9OvKCgCI89Prp2lqIrU1G
m9fDG8OYSKyx2OnFPzFnjwlMIybp99vPQ7aSvHDApw17zWSZCBje+LBRk8EzppNdiBeKf2T+AQB9
t0XN8CDMxivndgjWKgq8q6vXp81EGoiTkYc6Sk6AlKHCAV5hWdmbmDp5HMwJsBQa1RceAlKBzcaQ
z5fsYMI1Es3HEBl9dOOftOPaoI6/h9r8Ska829QrFBbwfwp+QSAneFIrbrqBWYVeQXtV3TdKIqKJ
RkTCDVus8dq89gig8NrGlOD4YAxv1/hkY9vTuVVCx0GIuURqYSbfQ6/vSvWMDe+J+7eMImyYutzL
we9TArdgbHP7lbBukA7evOO82h+u0udd0LCOi8i7l8PhC4kNNyeuhkFiZS7NLAdBuYvP3u252p9g
eir/rr/tntxRLDNDTqcIRBLQHQgOUXC4/0gv/fL/ACyar0wBBQ02amPB27s52mDlw5BeRCarKeEA
4j30CgWUK9zCvuqnVqCAdlenvWEFY2yXm+ADoJYiBbaQNP/Tv0DkfywuFthQ5kD6xRMf3gie02Cj
ETcveLmaLq/SCPNO+lgOhP/tzn95mYA8R8C/AKwPzKTEgU4DJj9FDqcOGQ51XDlsKcdK1JIqpq4p
/j4NwqyUQGjsDmHdbrGkr4J1UTNlGulPrdNYj8tKVeSIAob313cuGygo8YUZd4+5YL2IZ7tM3mKZ
g+6sy2lPGQNjIbYlVpHJFAVb4I6eaIB1iV36IwaDfysoYeRXkOTJ/iGXkHpvas3pz72af/HywWc2
ekQUCgQKt9uT8VnUl89VGEOEGMqDfQ412uQRYHw0PqxPIveROzlQrBYGgh0V5biPSxxFj+0JrWER
9nBlM9E/9jOMJpM0H6puvQvQS8svEPsY+ydT8qr7mcbIG5dJEOP0aBLRN3qfzllBlJUKFUtUazvs
mlmOkg4MTUQWJmGjz262FuOZptWytxWPe+5v6S2JiVfHLJgPf0JAA1HQyFgTkonkPgjrVztNaw+c
ld84zKrnWd42KHjhYtVRf+K6Mz5CW57vRbC0YDuORYTlhYtgX/IvqZe1j9/XDdgK4HY5NPi4EZqp
rvnXsNdSlVrXQ0jP8oKOSKMIHAqO3c/ubPny++ynCC1nEuEvszMh/LLkvQMTSQmznxKAawKiT+D3
GJgLnkqtGwNrSlY3Lt4+1Gc68VHR5bOX7kzhBCNbCxqw+uEGp1hM2ybcUUpkkLprIsYHJashjXCw
KGPK+DocaKSI2bzzes0jAh23fleeBAHAobnfBTOz3UQY4Up7b5cE+KqiVHlzegkIMMZ6eZMhHRqV
yx6HM7aj+QszTmGWlW1TvSJrwg2uz+f3EEh2vhGaasb1YHDEdUt2Mj/QrkozMTVVZHooreEftWlm
bhFLy9wUDsxguekSgQ1uQ4fQAueGcWowzs+s6IJFnVjDjCP7TG0B2zewF5bgrEFW3CEcQhgyOH1A
3RmnR2A5Cp8mCjysh72oyGgaMTW1fr2JOGER3ZgZQwKoya71vzPCMei5qw/P2v+nQ0Iv5FCBW/J3
ElyXF9FFGUVSOj12lmEePyYyM73/4skBEPwqdJ9SHPkoHvQjyGhS69CuxEb3hkKZ/x9WpetyZWhV
d/aSv+40u+scrupcvTucVQNUWGeWipTEjYmbNXah6t8864jDio7BGnJ9lXYbn+7iK6i1twOKFyY+
dB9mzEUN46MR29iwgsmDXh9sNsNfavtS+SKQW6uwDpv5+WESVd11Yvm99bpEiu9Okk7vFigssb+m
rUYXGoYdnR2Ph/RzR8Z+zbm6gnoENGmJYNRK23IdUlxKEHomIVw+//a5IYVplfvDuluzs30hyXB7
fB8VbwBThZTyNfXRXcN/pcDqFXt3Nu7CAR6lNNPC/R6fYF+raYpOblTXLTaePjAkkB+bBIt576o+
vEScJL2+9/RANpckL/WWl9zTygfzww9LsEE7+2CmT7eY7rGauPtvSyDUdOYSQmmEF73zcj8hzQZr
oa7dw2jjE/6CAimAdeZXs0eIUcaW0oHqMX17Q8oNLWjf8z0pFezZBAS8kdI6uN5xy/DX/dZX8JCh
xH4fvhPf5BO1EitACMP7DZIMIFIiXExYkPR1M+sG/YHYZ/FTyx/CTqLc6HJca/ciTMm1jgH2mKEO
eoUWrN3AAB5mcdwuc9vTaUC19i0342WKdDwGgkfUpWfONx3BvO5BbTgd9wy4c4sntTvgie7LyRv3
9nd07pP+T2PkiV1w4ZxDnhUCrPDxUHjxNRUZC5g1XOIvMGGkPhZSmTY5fz1Cbnix+2niQz5uSU9i
0hl8FTUKRz7CRfoop8Iz9MxIGJUhcKkwgSKJwwu/+AtdUbZ0OuKAO/6aJKxZRlDMeALYUiSMgba2
71RZ6OhjmOucI4ArX9OEpmkj87vURV7V4qqWqep2sLjsG8b2/gUOwmM7b0AtBzwiw9BfHI1hXiRL
kyP6eJXsEdj6HGWHvgvMBbFaBnqBGdKA5m7oCdsHFdt6DmZSYsv1nweuuOnXjjDqIUehQX1UQa7z
toR3/XopibQuu9VJkZcoSdDabm5HpRPXs/P/WpFi0pYsZvlTy6MfU9sSwMuK5Sf/UKHmn1+HveOG
znx/sqD2rkeXmfErqicfOKqA+7Jmpi5xcT8/wV+Cyl/gjbnGF7IuI7bpsaMTaKzqcg7Qv1F7Tbme
V2Xxb6zlPVHX8Cm/lrr2VAEKEH9+q8rDj3ST5TVcbIuLPfYjwMErcybhsdoYx9hW3zThgkh/tXOe
U0poBXKWV649OmcFyRrY1IuZVhef3tyNsivnOrtkVMjhy4P2E4dTuKEfxk3yo5ChUfIyWQX68S8H
qCGotL0etznVVGiVHT8wI3nnrdZWykqF2tw69stbsdbnZTv5mhyO6aC12bUyQROgouH3hgSrcZSv
lhSU72IFsWlv3lTtkJkVn0/hwgXKoubC/AjRM9b+Whr9b65IyYpWdtiGD5yTO/oKsPROP2ElNEN0
401bvigoBQuC7UhRju6bOk9GwfJTEi6R3tJ8k8t1P2zR9ptU6Jgx6iZ6ONoCOzEem0zWQwEw4H21
XyNm21sVlyf343HtkKuFCwxb2XBoD9Ul4W9rOWxVtSqLTPv31b2hdBayEb9z86em9nlUB+iRL51k
y1wL+oSkdAcD4YIbYeGgI0ZMLJQaU4REipcBif3MLj2mYSkgHcEbcHwg+gc6Y8gyVDTBanmiCdpu
WIFIKk1PcYVNz/Y0t9a0W7aUp000o85LsusLkrfDtdGfJpL0/Y/FSfFflIi/98tDoBUW5XhpxlNi
LrBGb/uTpKqrA3afqI5eVJPXdWyc4Y8l6XjP07uT2acm5wKT2VJH8nmJPttxHecGD5JA20U4vLK9
vmARNqqWOP/RelUGsASMJFl3npZrvgRHKkiT0tlZec7CBvtb8mJqCeYTODIgQ6XjThJN3UCo0xUR
mMH1evMlVCPo09ctsvhMjCJbfqDTUDrZLLi7GWnQ8NWF9BRwLL1Yi+VsYWCVAG7/12VmKoH9gu3g
nwRRONOak97IoPvBhdHmDEJz2E5d61sjwvwrdc9A/ZR/zEYgeQs2YH7pgYqxqzZhjonpf7syHIq8
lcA9/0YX1R5/7YJmau6lj9BaUWNqaMvmMhS7RvpWEKTWSM+OVyxEvsh2P32X1a3ZdM1ag5HN6W3f
hhcmvIrIAkP9+dXWsZ1oaLW3dwXvmkK49DPeScXN8cgeal/dtKXdn97NGBYV1kBuEPu8ae60IAn6
3ClqTslWjUiAlC6xTLnCJndRisP+NfKc5g3oYXsq31XFMTEGEQ/e5EqvOgDs2MuxyJ4CcLS0dYRc
fLO5F9tKHJDTQA6v2D/GgjTkr/EtAURwPKb+wTcxlQEVTzaCUYGgkjINlr6MKOSXedM3aSBxo/V5
DrX5L7ZzSqVhCgRWxA9WoGoTZT+FTu2wMayKWOf/7kFIPXZmnZEvcwpVnINWvec3xI9/Vuv8TZuO
ytvbSi3poWNUWmNS3zJuBPJoxmfnqgjURTBCYkwvbMKNLGQuEdPFgD8X5eGmRrkboKlUr1kj3h0U
SdayYr9mI+NdYFP4GlyekEvn9PpsuoR0ejcADsCL7glz0q0jmhtNqcX8uV+JBW6I46fo77RFfnQe
ZjjT1ZIgw3Mfd7xLvGx0oFArboNV9VnQLek35rmkWPV4PJ/3BzHzdkc8XOHmZWrMq+Iehoa2cAP2
nYNCLvE+WA/BtHiNjkHrxV60EhxG5yhQQk9p7G45boK97GO1Uw+IrahSmrnPh4UrTF2yTzfWAjWu
bDTfvPaH1nDpiC0OnUldtzyeN6ghAYp4puOrnjgmnQgcvQQRJX6oyZem/ap3lXAI/03PN+Mf2kSY
fUs8YTT9KyRoFHzdQTOfuR7dB3aeMXBjbiJUxI3Mt1Za3YKieBwp2rtRtLGdseTHJfmnvQgbvofi
x7W5LSJDPxW59wwwtwkC3cT0nBTTdNvq6JOfat+MaWG5jtaFkJ3soJYvGVtuMHeUvzv/9TupgCoU
2e8jtM+kSRqaIhaZLWXTvxhGBB8hnsITPyrYTZAu+Szszi2Ona4+cIgJbIZh/lqeG1xh+84uCMJ9
7MlvVlz0GMlqVH5CtFYehw70mdYt22nO50kuLKN37Zxy1Zin0Skb1f91vh5dakX5xEw8gd3V6tfU
UQIa4JdZ2P8LzCNMaMvuXyJ024drI5ZyE8SaVgSgMWRHWsXVP4GehnbwN0yN0Pyl4PAlXmdgpkiT
cd+ElSv4lsLPKk3/OZjS/jCZVyhPoPBWLut+qrbmt1a01bufzA+znJHbxlcR8PI5n8chgfTrNYIt
CUmMoi9zM+6s82pky+vGDQLfMXjTXCPqCKNa69ZrScgOkU7+T4CbYIe0O0XDrD744Sr5E5a0yvQb
GY4MNvwdGBH17lNjMlC/Z8F57Y8N09i/dpiWOyXRB5VYVX+lB6Jdxu9x0MkZqHOxUmM6fKP5dsAN
bhIcJ/mNJjWbCd3E4ZwdX6Y2lmELYhtH62jn3AP+FlMdXldsXACfZ//n7ZXx96yw0ZwMgVg7W7fE
VLPpLSdKujy41nT0+U5Vst7lw5xWrsKYQIirYLE1jUvSipO8G3hNKcb/h1Waw+lqP/UHRG6aQl3k
2x8uLdl02nk9F+IstCwj36TYKTQIbSvLfp1X+B6jbk+98Yx6Wl3qfLJZu54cpQrNmDWLp8A0xyOp
e2gBadbYW7GiU52wi5Vi1yDJ1eO2OvezSi++McrERLgZueih4eUdnz1cd7xmVFj67LXdxzCbyIbl
zauVWkrVixmoOBqEJp4MLLAPQE/AB9AdXc5nnRTjV3WEEiMBGYKKjEqGi4ASovdX6FjJQzLGZxf7
UDhulaVXsDSJXm/Omgr4rGrDPcMxAnZrCOwrjK1tzFspRQBsaj6QfcKjCvhZSQcNkz+eqMswVlsW
BNyrTeOolL1Y4zB7fvzk+VJNCxrNJdi3nTQbigvZk3sEjeMf4KWPeQiH4OkuzrosEMeWPqTMlbkJ
ChNkUf+OdVEfKShgt2PunX/7njU3jrYJf4kYpKacFcO2B5rww8SiNHsbarvogWrLVfgWbHf1KO6K
feYceGcuXvz7FiZDWMpZUTPBfMDrmYAPOFy5Jte8lZjTDTuwakHUcxeteConv3CsWtAXouSUATwn
v2qXnsIH2OTObazrDhOuQEUfPsAyyyIHafSKpwPLvGEMy7tF2LTR6iVJphgmRq/yLi4OHgfnvrqs
MAQ+nXvv1kahzyO6YTvRfCQ0J7VgxrZyVYAQUb7ow8Zhl1P0l+GEpUxFgrjiT9mSXWAkHj/1CE1C
aplv4B06xbcGKWjN3IiS0irGB6vOvjhZspNox2qPs95bRw/8kENnDF/ZaZOjsmOlhI0LTuYa0Dj1
v1RqMj4eaeQgsWB5wcpZ/uExsvYThnP+HNGAi6NjoJIkPI3FUO1Qj3j6CFzyb26s3BTAMDuPpGbH
GH5WCsLG3v+3C36fhYhTiqylhkBHBFQeDI4y0Lpo4VtqmsTN0o4dWekO9vhElnECMZqh96465xQa
JRUdrqwO+7RLF0BzUYNgF6KdS3mLmT3isquzEql50AAOSg/3XF5xfVGYubHicZjCdW2dy0FB5P4r
f1Z4jANd+Or/lkKg3jVzqhbVH2CkSbms5Q6wb9Cd/VMoXBN6aw/Xa4i3DxgBkxXBTzbujfbGgLkv
sGagQ5YYLgBTR6jkTmHs2Q/KaqYwC3yKV9C3Z41j6zjLaR9iqHPILUYF2lJfd8IslNJ0uF1eG/5D
jE8ppXULsOGXQOuon53IhMWVMvP3lltnflXhW0DxrEpmP5nSrs3noC8B3cyf0GHH+QS2hrFDC3eC
grjoJEy1Ao1bEc1EL9mo3Lk/t6EhPPz9CRqfT+QGUfTi+QwNi+NuAJLpakwV4jRnNA+yfPEiQ4/4
ojFy4Atl8esbYbIg268o2I+TJodUJ0hMbsUgikQwKCLN4pxE4FvrknsxnXIdxxqflOeFdzYDsNTU
Sscy5jeuvyI2Sjyuimey2VHGXhCbsQiQHQGGhZuncIJ7+kO2SkAiW/J3VKoNf+XHH1NUGAE32kx2
ZBQ3nCuc42OSoLvjLQ1JsN18wHYPNaFOjfh1STJEkV41O8S8z+D3jv5ovpd1XFoMjtZ484+ieR27
XelDarMXN9nlxhRVJgqDalWn7E7982502ucSZ2RjAesaIFUTpJ1r9FOjsWVmSqqQnRg7kCGNr0Nt
eJeRURi4Ly32bNd1JxT6tzChy4IAOT9lZE3d8ULUY66DVJ3nJk/w8FTsCyq2jwdRgkKU3u5zuERE
DyA44/6too4q64lVX/65MUu4CeGcB67GgfmA3krZdteIUFzhkKqNn7GEzIiD+tdqSSVON9fJTmWf
9PKXeSIMfFV1Metfy4Sl+/Z+OW3DEAm1tAJsF/q6+h6ilIW/zyOz8yuJhZ9p42gpu6jLxWsgctQA
7yW8uBwlrL2WjsF2Gba2kOZ80iGBj7FpXzDIUC1PKUqVmv+QeGr3VTRQMNYBojOLL1QwFeOljYVZ
1X3ZT5+ydtXmCTNuCuXKBuEcFwh9Ystnsae0fJLmNhe9W/vLIpwKh6kNUaJsokAH87nJrQGpR+di
bypNYVA+jztlOZW2zKi3ZI8W8bB2SitmN8uN9OHuqhyXQ1s8XpSirptT3MLt8OHtRlyTuwwR0lw/
hMr4zL8jA0zYJFRN8gHE05wT4uTMYJlRmmKRGWCbW2BI5jfgrAliF4Nlw+jIjB06RAszomU+GbHb
HoCiaqMAlzsu5pBotO+u55hgMZU06ln+hxh/rz06P85yOYSgHFS7QK6EjsRGhX+nP9jD8pO0mGTu
KK6vpyG7myLvT/ki2iKBhaiZRgN1eMKQoIAi6WmiJnj6NLv8qd+ESvPunOh/Zj1tV2B8jzDdvi3u
qwZ0+DDXPI7GWeuGEMRjWgr/OOlSkNfYPWaX7cHMEZ8dWq6U26EzCRtrJHhdU7C70NZhzoPKMYTp
72c4JEOy9eld+8VLOQfaz3XTV4+5svz1ts0EJVcmUSUlY4Sg4yKLDhB6fG5UE7+sWQnC2JwflbJC
U1dlyT4N1PWTzwQd6a7Nqa+sSjk9RcEv0xbolHJeBbuMzfa5GnJoqrm51z8Y9a6WW4Yf3ZZ9E5fQ
vNxNMmbIytHgHtO8p3kyGM5+94ph4GfysjssUzLsi+fUWv99FGjrDBHjxhtABCm2NUSJxcrbEnco
9QMGR0/ISgrhhDkljlR9wijx84/ijZUE1x5fmsmONUcjmjHBMTn2tTwE7e+1Z0INEnbzxvic2ztI
n63RQBQuVrcpz9oQDNmRB3kjn5Rzlayr6KHU8+04pxilM+5gqkzgRpzl0IRv9ZOQVhvHI8ePNV8W
+Cg9Od6ud9AfTIq5rllRRbAz8aQOF7u3pzqzgRE0Cm5+qEeruRzmtQHZCgLAm0GsCs+/oKdIK31Y
6D5UUffC2G1rTcd0WYbfxvtAka3jBMpl8oBaYTqHloV7MB3UBMKTIR+5vZ0yHekruN3JR2npsg6k
2Zt27URtTB/PvX2eDhFDqB3NIV2Ue3KoaJl0gNHRn18AvgLHc7dqTsVnTX+77WvL+dO0Aqbe7WgF
OkQOC6xEI8MZWtNtK5HZYfseUPSQzgLFk8d10PTOb06vD56fuCa82VcnmQRzmEzB9BocLSe8COKS
RU66r+EBX2soUNbTMe7+3zmdyCjCa6eOkA+usjjvWjY19Lq6PnNo8hii0oJEHYNy/X7I2uuqEax8
KQBfu0aX0p9CishJVJ2Mx4ei7qPMbIVDTRaoqRKzIdUmz8tK+I63h2wBVKJ7CCcw8g0FPSepNvL7
Bb3ortIDysmTFNg+f2YKDcWU3uM1eUxV8p48iGPMI/gxDEnGA2MhBU5MnyWKvWhl6BwyGCbHFD3B
3glj4Doa7MhoBYN/8VRMqWZk2bIoF70Qvgu191EEwVeeT2iTPt/cBnJltusbCzjI7Ts49wYjoxC+
eYbhF9DOz/ScZxe8kQpzLNiOvPC1cYGEfPpJwJbfZDpW9/bAJOGdpH4QlaNkxqiv6hqLjmWEq9C1
JTp/s3MCUPLEJpxxT+UdJyqhXGhkYTp/kI7Ibxs4FzuhJ7K7rUia/UFfnn7Se58ROk4ldAsF4mPR
dPtZ+Iu0gKoRfQYK/LlBGY2LxbvEufJwxh5QgNUTdz3VaFIxTpXLhXPnNE5wJYuPYTJc+xmaveOR
A2ULTJFVKleqeFUs9Ez1/kpYoVFsKT5bFqhjvwQXOsBJbA1gBLilfLknKhuXegs9ME8WkGFOw0IH
xUOANcZkBLQuAUz9HShWCtbxvNSVW9ODq3Q5ATAL/7advXSMOHBK8X1YdqyFbA77ChQ+qShBuN+Y
uuWTIpqX9pxKH1foF8y5dpCVMTtR0MamklkbXHilP0zPO4pF9KJ/+/RsdHqjmnRc5wk8xx+Ln521
2F1eLXs9X64L+1gI1lSuvVvt4IX2gTo/OEZeFHIf3BeNB1oU5TRsAxW70OhAIP/rMTfsy/br3C6L
T6e5tz9PAnuvzXRmB15hGd3mhRe/fuCXFgovF+9lBt59uQWBbVz/XWxESzQnPiKv4zCYpmK6LdUk
0p7XG7ym1puWIIrEby81rqUxypSjzkpHn99GKsZ7vVKiWMimDRRYlyuIwanEqQV95h7FvgEzNMbj
RSH+5X5crwXBPR2xUJ3HJQ/U9MQpPT5PB1W+maHJvXQGTIU3VT1hExZnCYaY5d+46KoB4DywgIQf
C4SE/CxaNR+3dpvTwT8MGA4MNHvjsZ+VHkTfiOWFyLAefJR3qe3AsXlU8/L0H+I1cFx7L07CPxNI
OA7iMSHOX1Gwlq3Fho1e9PxkLiebEtbPtae1y5r+zC4s49SmAVSr4we1JWEAkAO/MgkNcQlAKlbv
JZlH26h6IBBJtiBPqcti9Jqe3nDDOzFzQf/CCUIdx1q4scLV0KHPL/Ve7DDI3KdahkXo7rapHJng
aUbPEOog/BVsktU/BPOv3M3ImW5/vHKC4FP6uNqp4+LQk2ZwMC3oDynuWLIr8cBSpZl3MbT3hv5q
ufv0c+hJHuFU1AGJx81DAInQ/xNIgje9lDlfIQRufHCY8+AEW3+h9PsiHBo/daVvkXvul9le8imw
RH9ilXvGUndIiwy9XX7v9v5RMGK5GxWRxkWImJhyjmhXDcYzpf+KRaoUqQRd2QM2sHoZN+Dic51k
IdOBae+rpgk/TbXGcK3+uNZ8+RJZf+LcVm/9BaOXs2qNLI9k/Xdr7M+7XeFq7sfaC0lRh23IGiOB
PMyGIS51mm4XnudeSotOJsCPW5x28y3CE/M95sSmS1hy1royfaYAnggdEKPUundZKaocaTjlkyeO
8QQqBVasos6o2sWxzVQV9unx2ZBm2n5DdC+xQ7PxQgLrr+eK2Vd2LEOpjDEWBxJanMqAKRkWQqEu
XrxYHeRNUkDN5RwadAASjXESXv4TeciQNBJH+YjaCRC0wH4QrcJ6eks7hubR4f0IvEDcb2dISp00
bINNUuxmBKl9CUM+NP2OazlOIvF+owfbE7jbzP63dMShuwTfPsLpgE2BFueuVpqcI2VWVuet1MwM
LnbJar/2rkE0RqD/WpypeCGs/fDU8fZePqgRB4RLFUKydn/Aawy4CZJ79S1ZdlJSzgafeqRDOCxL
lSu0MOQGluPRgiJY9VJfd5koT/cto1jr2vhR6SW+H+Wlj+Hk0DT4zpiGPTAjQh96uTF4RE/mcA0X
9LrQHyTUVqPI0BH+Tcy/UMVx8qX7i7QBOvzq0OxbudqsKBbSOCECNTBr07bygaXhQDa7ciOyRenA
qYWZx0AepeG0ExBhr0hiq3EsQTV6RekA/+94yVRamMlvskSUPxrxI/zSP2gOk44rNKbYG3ATUYEp
d3B1JqQK0DesqxQsrgnT2mAg+b3xJpG1FHWAP31/gaQnJ9I8EHoVHbrIQgN3QK6Ay9C3q8v0DXtR
+K0vxbFbWmmK9WihZFadFAWd2lJ08fcKn/mHQF3K4Pi+3xzbk8v0AA9pThHhYcfvNcbHs31ZgyHv
H0502NAg4KPptvNZhWPDn6MUYZ0rLzHm07TihPa9R8bcRlBTMEE91yE+9GjLcM6PcNEUU6Yu4APO
3W06wyTtYH9BoJCju4E64GwsbEaT3u4C90F8uLWdi1QNXVWTlVk2pb3HPWj0mJ/OiKU84VN6YOg6
nywXyDWVxm5HWaUIOPl1KYvDKgMHGkbkOHqZKEteCcg+uUY6ljdw4Hl7w2UnqNIvayzEhCKNLcgk
BFsxo2+oQwKFhEYr/Pz6LaiIrUXEV+Z04/WR/N8YbC33rlkgPrT06I8w0+YTqrjCM6x4lL+LaHjf
G2nq2TgWoNlw/9dOWMIwDS0cxN1fqtLSZIdvMpV/woRjKJTHrEtn5cXBSY1qYgraoITZN2QGP2x0
e+D0c+cSZ3A6hzGSNsfs8dIn+gjPqsOL45daWLjXppO1w3mW/hz1RIBn0cfV46ridz6sy64dZ+5g
VhLyaxHX3ujRhRMjYKebYAmWzCcrp87tM7YSkepy301l8z8gX0EcSje5JS21djLevV+2pryqgWyd
Mj9p1+2ZLgsTwXlKv4ELgUskb0e5Kto0k0bZPh5MWhB+4t4ZlKw7vRLsjYbgXkZNCsuH0IlMUXlR
mbpSmxlsW99GHrl3M8GZR9O/V5tJzlJFfRV1IKgCIH89btCQVUn1hp6iNqFwUKxBog2lX/0ClaT9
NF4jA7imsqGk9rwN8LVtCQS1J3W290iyyWVPatIZVpZODgvoPCml+A3cvfPrMs90yLjDTYYQf4+4
gxQU+StgoZyGDFtw652bfHq0uiko/HY40jQAiZKBT+/7cs9HUKL/wWV+q6U4IVVG2VUIgl7JGmax
jwdtKKBxj/o3Fth2/9RGuLON5txtkVzEdLAeEKTWlGet7pNkUouREzSat2ZXWERRdogi1bwmbrpw
os0JeAw5Y/G5BXm2x0ccogBuMvyUPHlYQOAPZ44mALJfaXTBO6mnfMq8KNRAXk+A6pqlAsdns7uV
beY+mRsoLL59eAqANiB6TVzmAFq3atOPF6zAkegL9iU/IIecErAmr5i+eadNLAQWlpLr/z4TGePo
C0fdW9w6EVkqSDyenxTI9nDO34PjBUEbafUlNg2QrlBa0gmpWEqD757dRoMmwgGI8kYWK+/PT7Er
NrWPglayA6sWkRd/lzzjWNPAjoxs3LEq9YcHu2cppa4ecngX4uRR/pbElB8Ztahyfh3tN8xgUSoO
SzjfELe2N+CU/SSzehVYhdNuUMY0JzCGE5sBynBfzSGjPP3AWrC+FJbW2DD/DF9Mpcjdo0W074le
4SM4TsePXU/hPkfCWpoe+Th6r0TxTNkkjU9A2WDOFAWS/MFwUjmqDxbEreP9W6CDaKQL32tOPivz
eGQLa1ctRNPAvZPg/Mu8F1tegIrmiUGZkuWE/cTzojykMtKENlj0n1bFsW0lrfqsdKaIX6LKpcxX
WqOGngEhSNvb1JvsZGr5erxhQEVADLfGLnza/coadw8eReIKHVUXgg0RIhnwgdDU3UJ6yCYLyBUf
DmFcVj5yzImIFrSIR2Ka+9dppg0qCkoDq/8925Ps2l6NRv/E1J9xl5cIqSCCZGJVHoOWTHguW88E
GYvtbOka7f853E9/rBTdaxMDcywsglpZKHp1gSoyoJcPQfE3RmzS6hNN8RiAZJQmYZ0CbeicXEYg
IkfuTgNAW70dTeb09DG9YsAyggJ0+DPtRQA0MrD/2nXD8OO3782uz6z7xYXIE6qLnS4QJUaF4uxA
wM6qLYIU0JCgpclNDNw+meKB2euLfdLZxlh0bUn9C54Y5KZIbzF6VGpssYdB2xhamCkQkdUX1JHK
6Y+/BHKaSehlHBQCQL63jN3lCaZJ4J/MYViSqpasSz6MP6haVlDJ2jNrcYrI+J2F/CGQV6RvqaVq
LlvBNhWl90AiCF3d+uCbG0PhYbr+5XsMhYzpdDzuPAzHYLTNAXg6CeoyMCjzfrIL+gtuqp9xc6HD
C4MNNgJlRqjlcV4ywwJQUZ8RjUwBX3KZSSTEagBAhlyq4PE2ZbhTj9xpESpAdiUVp/ullQ5E1XnC
D3RbR64mcFnzpwUObtkxZwE9zNjPbQDiG2Qzk+7nMfEuFDaIaQUbd1zFpwm+3oisUMHpRgWHjTAw
of3cHMRHZDeczhirdyDKtOgH+7AU3q30BUZC3g8A6F6MI6SKlzAvzpPDOTDqAOt/dSDQcOaaLc94
YnXnPo2tbgc3Klmn9iEtiYBbXLvxwFeK7eA6wVpA3AT8APhfHHsfXpMWrDHRhaxZkhVCs9C0ZzTh
HkPC19VHdJuo39HlsKzbcitcna1L/5EyiY+DtWvWHF/oN131gR9aw8ASUyvjbNweJZnItcMDZRa1
wwAzn3J2k2XHDqybR8myYu1aDKIan5Ikn0dSagg67NrC6Lk33H+1x0EKdTvqPxEKuEti5svSrrkv
3JsEjmfB5iHclH7eBQ8exAp/jDMpFdYRaIkxDq+Ibo7XnOBMTVnXOcenOFkm6CgfRFsNDUMbg3T2
UOLz1bUqlGZ21Y1Un/AVmKkYkI1igTHutTfaLdd8i3FEsDlYcBa5iUk3fzOyK+afEoX+9sBfGyGT
6kJhfoHWDzuAQ5f2IcVchqBksenf03cFYsU1v8wsSo306rniq/d28z6Q35So4Mq5PmX97F4m+2Iq
vT0kuXC1m871AfDrVGfS6F+Aj6BG8HbuhUZx7+4PG6SuozCrXWT72DCP9uo6i2nbEebQQqnvvHdi
ZKCajIakdAfuQMYJt9YEqkz3QeLwvSRiBAkqvBOcTxjkc3ma/rF7vbT5idtBcUrCxVF8Pqvycqy3
IIG/7gSjvDQOn2Rr6Q/PfxAOKaqD3ohq7DVw7gPsjyjQVgGYaK04M0HMR2BAJygQubC5+pZIAUHo
3jm6w4lQPPOSVPt8MOlu7Y6QN3xRWxwssfZ4oyDUSrZ3P31/2DQ3sLRYldcKVz3yIeieZ1u2bCPq
GViLrw4WEeWPN1wgKvgL7fsCI/0WLXj+jDfirTuZGIkJkE2IBoG+oOjqvlF4Lth2M9ppbmjVwsPK
SAyfUDZ1+yWiMY59xHfWNEF1ZYpkE3I5SApJm761w9nVHVVdIdvP4YDsQvGPgfyfuu09y6NKZBjJ
8asymJMAtskWn87VZyust22yQLFQ9NNy67jnXYjRZS4dwhIoB3jDZ1k46FE/8/qro4lXy9nyqUKw
yXLVWI+2eZm3eyYqZag8XKozbK81oxOy09UCjyErDytQRfG5jL7wm1bKCecx9VGqA2kMJpwNc+GR
sx8FMp0e1OCl/EtiTu7Gz/3ydSfvwsxCA/W/wsHxJRxM+x4kj+6qMZmmAecJW795eDEnt2CvJqNu
pnE0vo16+jwbZ9KlzWLGMlM3nCln1hPcms2NYiI7s0w9dNxwtiMDU+S1Q4qtRozHJSN4ovua9tk+
xpW9Yk8HsV6wy4ydr7D4b5SuaKfGB9Sv3mT+qVCwZyYfQDpUxbIrQGPgM8l/msdpBxW7oJ+xbley
kGzXxRr7kLtn//gPCt4fMV/fCd0U+xq3KHK4jvm6afp8fz8tGQcHrQkkwdBFtqIbfu9c/X/gvQTF
B0fxmcvFJbZwihSFl2RAmjUyfLViH4XGP0U/zrMKXibsyDmc+rEPq/uTFhxKUpM/jPKaE/TM/79C
tov1hGV7XHdDOYSvFg/l5SthCUWEJWq5POAc20wyv/+mmP1Te136k3DWoLhuaAgOrTz4fbbhukPD
YkM4ZrLegvhqQ2Uoa+v+ZWWiTKXC1FZtaMo5LnFd+orgmrPkr36AwJZWRfwEZNnMnI89+UqQtmG6
jprVLcDI6Td/MDDDebbH35rZx5eNtY2G6tmKpSn+psfMqyn3YElmLuYoKyUZ0XpWGxrJwZJv/TEk
vcZQ12BOGoy89bhOUHfForj2L8wtDHh+WxeHlJPTk1+GVBw1gyLUyqj8udnITl66G6LrexP0FkES
9+O8KQgzx082kRR2sK1IM68kolNYLM1pMO/vTxcXzXuLecqJB0df6IwlFTldJbq6pOmjeXIPChQZ
0p+cfc29Mq7YMIeAgIWOevKQSOC/+hUy/MqEWJXnjOGNiUIs+aDL2FTVQyW6XyI5DOsC7Q9RDRLT
ZTAm/JD3QduIWZaHRLETZRGDJLMk/vJgEK33bGMjZSYt/0ES6jnx1Ys4GcZB9GFzFtzl3pUsm5GM
y5QZs20FL7lfNTZzewXLQ6dPsmQcccywMlGep6d/EhV7LvX1VfBnDfjiN4UAaCjJagNGxVgeYtdv
A4izCtJTmZ//2MjHwG0TS8UG/3dT6hVAvMSyrO1PK5POyjns2ppSjlZmYwT3vFRNot6O8bWlKz7q
ODp7FHEC9XuFhhPCwojPqSnW0PCTn/t0OJMrry1b1wem5C+RqTSgW+1BG8PDykimHq1WOi+/viyW
/cL+5cfO44RGddNsGRvz1LR0XpvYkI5ElZP/6NHu2OEqKke1Jh9ryNwbeMUK6jKTcNHL2Z0OIvAV
lz/sC9BzOVOaH2qtirkktA6xXC8NNABkiCuwaJ5iIKBGPL36g7ihZpP5nOZACmyzF2fBiGBhI35d
vrypGDZwcxweQWEOmRYeU01FDvAMAEVO5kvROqFrmZePFKV+lFLxsG4RhXEZN40fb7sfmITXPTIm
bgDXhnjIUfEcMBrN2wMUbVIOSIhq2NCwwfvGf7XW3CV+6ttsjyTf/5+IGUBstZeM0s5a+hQewcde
6ijpGG8cOXvFozActr3T6mwdv80/NnNenyWvkIbpt/PEa7IMqwL4nr0XCX7pEet1E5DHf4g5k71L
N/CbYz6I50Wexk0yB7bukZnNUoxVQZsZvcfo788jpFrzu9caOM0dMyfqjsoP495n0B0Twht8fCMC
P7hdauyHi6VM8Q8cp1CL3xIFC4TZy2JTwJJa2C1LSMlUhm5nfebR8yX5B1nCs3ft360RdtvHEsBq
EbRT9LL7B1MzwI5YeubR41Z7AkNH6CD6jqrbhr+wIfq2QrPwNIVIrKED03FDvbSOn9TUdq7cF1kf
uTYbAwPQy+NobEps+id9lhz1lM2PXjCBiwvQt472BRPJBTxNCN6j1R8Oaw0imKzkh+JuCnF5zshm
4t+pQ56wC5vKZKg/OZYuIWG8/q4UEnrLBzNZZ+7KniaN9P2uwh+yebaryjzvLvsKBRiROPCsSAEl
v7s7TWI24FX0kz7AK3zZSImVBdJIfxNSA1BYPaOGAviqmhNl7NbPgfM7lDhvyaUDjua5fuQnrWJm
s3Iq3v2ABtxyi+uON6aH92olDDCyWjrrAsCA+/olyN8OG7Teweuamdk6kJRF11WeW4KkBLSTIeVZ
Vh6IEBgssovilEpkLFmmzabu5XT4aTxvhsjoue6u5RdfwH8tonFsdOh5HMUTid9oS2BToLyPqSSl
+A9ds6JvNPTBsCwyFrBraRHEkC02FeUHf3W2z5LNGcKBUKqEqFHAKCFJ7NlaWUNR187mtVa6L06I
KdEj2ZYtvNm8QfRXFoij//LsapGAWuMa+YcYmIQH13GNRSRqFD3W4mR0W/7qJBKMnfUYCWPEQAMM
6yHq2eWEJwejOdOjNSuU2KB/ygmYm+q7UUCpsa8ADfs9FOXWGWoRIOI+HTcOgu1XQZrRK9XAYPOI
rihZCFTBMiqeOhPon7iKHOl63RXQb9fE8JnJN28Lo8IkCGELlbhz2NSbkqQaSYCJ1sQbJZv69MvV
h3PWhOLbnFEBbybiy86WeRfCgJG+lkG7/614D5FX02Mb+dwCC/NAunoWg+xoQJ+cpMIWYkNp8MFW
OZf4FXLuiC39u/uqO/dNT+17hSFQ6Q1bsdFvAh7/udomIhy55WUdoOUxFnGEhq1t+RhWopOK6rAv
izns3pHCpUC4eKK1d2ibPHr4w04yTQo72jWA7qcZxOKmfpykAM9KNjZT23aDAH6n89514/taNLBu
xG+vssn3mh6wPOygYz+ybwHsUnJ6MmMFv8jLhYh/K4+I4eLNQAvcd6ziel6Sczq3QXedFkEmWhgY
GncYBK38LliXH5J17JEaYNADtiTReF3YGpJjF6lLgyQqM/6SmD0n/V6qI1CckBZ2757CE5oFIx7E
vsYwe9wFGt3zfmx0razOnspvDOWioAUYAXm24V+PKjTvzr9yvAoj3Qb9Kj0JSuaU9izh6xWzLbp5
0fdWKCayAxTkEQQdTi1d7fyTXN5QkXs2XG/LOEzpZZcNr78gnK8YYA8TnI34vZWjqpGYsopGowwP
wpWcwHcBTn6trvq3VPrnOYjwfdoBeVl4+UGpynkBTDAAWKD31SbBzwe7W5chclV3EboJXvXk5H1i
ZIwCgJSMNa0QRI5IK98JqmfTm+TaZR2X1hSYeAOpwCJL13sRdAdPsenw/3dlgbJUFTkBFcPB1LAC
8WgjzONQouLEWqwC0W81hPax1yoxq9ntZhYosj2tYd6PbrK/7QsctNFw08bLk+QmiD2gbdAI+odi
ltFvbEIUOrJjfXy4RwYBNN+GAZhOyzemY2deQhR5JFhBicCjEjgO6ZwUBGNgDxa0YqwzDUlOaEhq
lB/Tzx3tBOAS/pI6QHZg8z4e7fPh+z37/nD+4Ls5Lq7LuI7zIFkpiJZbu21N9FDAfhbdjQOPk2S8
fQk9ZA/jyT72T7DZUgZ+4m/eoa1Yw3iMN1g1ANwnNkbuFhRieRZCJWtqn/jA5CegDmU5Z4pdjV4C
Ph5DEUWoJUiNd14pds9E+K5if2/dgY4bhpilKzcwKKC2WShSh3F9xASPkMLNb5/ucAhKfgNIMGwA
8Uw3l2+Upx1v4ywHWnWm5HWLJ1Fn24qoDdJruiIHnicnYEWpntl8a1lGqdD+EJpWGlbmFrFxNBu9
9AMKFxSoVurbPNWtYYPq00s+Cb284NPtxhQiOdW4WD//5lk3mzfJew3iSafq5RDoENitaq/N8i4x
f8nghiBbGQUAmXTpQ4+LEKjFSmg6SsU4RogUZj/rrZ2jjNe2mnQOxo/xiy25lW6jfqyxu1JDYwgL
g+sgi+vkLu8iAr9SfcgvaCEV/wg2UPwuVKuOLdDItqv99f/+wKwNiYoHfCCxZwrgO+Hce87d4VIK
OJqKYUySHaPjFymNxgFFzGERAcpp+btkBbtnc3UDaYAZxNhCl90Ch0dhaW61AZ7yWGIMXlehmx1u
okJIoMjIMza2Yl2s9dGuIB4y0DyDep8Uh1by5JkcEhDZrgarKvp95O5jfAPmXmHcKPWFxRhPSZqW
p4SBS04L5zPIe/sg/vN3qiWpErxw65n1ZpooYLQQeF2hrFz2jzb9YUG8vxBV8kIg09EGYJrlv0gp
rc8PeyH9Gt3ped4Wuq0i64fJvOEe51M8TMK11K7ylh3W9zj+OmxDKaNnbPviwTbOCAPHjD07IzzI
UJm4ch8UrE6cpvECOMKvhaL38rKXc2YGSqCPQ5RcVPSDytp/zNxgU9P8KgCkCR3eyEjCrT4oeTJH
VqEOycISQY7Vue2RgyVOffY71LAbTWtCfTbkhYptACP7Wp996jxdoI+k+c5PxWJ2bF6E32/vuV8Y
YMMHSAPNDVBy25jYowHddactb00kZZNAz6iOeWk25eglIXIBtkeowgyWOmcmE/k8b1usi0gElBIF
ENdu87kE2wyjmj1mKRgklftLrZHVpxLVTQgoIlHTfLqJT7tG1MDWu2UjZ3LDAKouxz5i4jZ27UI9
CD3TKA+7rfpej0eqbZ7rZoWoiicod3FIpbFr5s9kQT8vbeLLbobc8x0HojAva4/hhn27TUiTwezI
s5zzIIe5xWjtOAGnsBw6pcCcHL4nSNJgHVBJgtMizBP8YGc1tX0ergWgfiR748NewtnJmX9MUgEn
Muh2MwmveWRqJhEIHokxUahEU/WAyjtQJ1CtRx9m/AJiN9Wk2hUJSZeMXN6U1TOK5fqyr+ZCICyz
9WuU1k3yumMwGlVTqJybxPrVnbOrZTi/uNoSSj/+yn7M6gzLglinjR81glfJpKri1aTfsl7Kh8jq
61jlKv8P1kRe9dpei//zbc/55Q9aKAW59eE9NzLBnJnSQQdVaAu8JB3Lxb6VM5ChkcZMY0u749+2
Ibwi78p/QtoxN8KFvRDdYGIolUR6fPrHRzycHpGNB6nJqpEkWMArReTu6WWkoWYfoGT1+WK9fvlX
3N+fLz77x4eA6aQEiiJZnl8uxkIAQUkRs+VjPsLwWpZgY465MCiQe0uIBhhQojsTMNXYroUmnevc
iJ10FmksAMBUqgVKeHjHpXgkzp7w4gLDJ98KCoeTgTG01okyxL3RE41Tad6G+s+YVZnBl/ak7Lam
OmgDsrSyr+kJhYtbFlEWZtDllazOnWSYAkJjjJQetreupb3gEBMlqkqEpwr/loDt4XIyoLAt+n/H
HUU5jVVVmEoM/+2AGHKKkDGM7du+ObPG1nlPRBZpatl59BINxwIVV1oOoGsTmnOe3+x9k374LIuc
FW7pqtaCG+xeRjAwpWcrFyDZ9U+DY+meo5RU1NalbMaMny40K1WPzjaqT7beFy6LwrdFa3CjxmYQ
2tGiiIYXB1S2EYoZY+/GrTxqBxFrBIh/BnneyKMaqvS/b+XeyReJbp6RNuitrBM/fg9AK7lxveGL
qPyb6uyAEYiWsD7pFXXEudgwzrUc4BJgfufJwUYZJuZl0hK3VhkoFaGGVP/yvCtLwljStUpgby7l
jcqWrsEBeVgs8OYLfUufZGgCZtdGwDuF5xmbag4LPH59d2BnUQJPcTN2rFaktpQb1CWzhcJeY10u
6ERvRbhlSG0pMl0UOO4G5AQ4A8366jOTvVxWuFxpUG2QHWnE17vIdyO7GWhFgklVpIUTtrPR0ThB
x7P8QXQE/8CwWhXP+ZafJBC+0e+rEjDyWoBeq97PNnE58VTv52/UH/csJXQmcB+jAorsrOAbL68f
03ybx1rZCMaYkH3Ybf0GF8nxUfYM8ZAHzTS0jRqBQfDOAbnjaHcZesb1dsitbvl1fVGk96eDbUR/
zAU6VWFhnzYruthOAiR7Z327wwYdVJ77qlf42Qkqkc5fRPFoULKJTg2/vyL2Hj086UFIiBkrSoJE
PXkLVYvle3BakpzNLr+JTtia9Y3gdOvDRw90hkgX4/SV95TMM7AjWX59OeOYDRmKBLyMWXEQ1X5H
wjebDSCmap94BVGrbwro1X6IY9dqu3ORrkSwaCPCr4pZKueCqP4p4rIPs4tG9PLtw6eMT9dTn2FK
O7k3d+9NiCJQbA+qk1icHPu9gl46QTHfjn+cfyJemswstVbWh7bo5eoqxmIPz0fkxNu4ojL2C6xm
eePDm1MFqFiAdddgT1OSfDwzj9q0y6VTlmywv+t3Qi68PNNAWDmlZdNv2yEXDOWoWDCxWE7KEdgp
twu67IoxkFkZMl7HKDyGheuy2121y/BATZVmkLtYs1YYnLC3pm/yxe2cZ63gSzZv3KJeNENU1Xaf
U6xMAWYcNkoaoLfhqT8Z4J4DwvTalItaodTcs8OTWW6tK/j/JDJJOkx6gpKrvSyYx2hEpJ9tySY/
iPZmD6LfdjbKc443XYuino2zIBMNMpHKAXYUX1iSa7Xqkm1189BfIlWSAYafxY//uVwolvQVMH76
HXRCFq4RZHuwjFq05iL8KYKNJaY68dFGBV5dnLDLLPyiKRVSjBqvbJ0SY5T1NmKgRWF5C1xM0qt5
ziywhKN6mK5aITx3LWt8vh3G8YN3vj8GiX0NBPf++I7AqCd8dUdYm0w9HB9yRfDn2gQB25+48/tQ
fJPSI4DHF40Yf1FPmEUM29s01P3oxGR96qoNBBw61rRk2OeEkB/v88fCWXIa206GlH18TdNGU2Y/
nnpoZ7zgi4YNS7incyLsOUOPvv3hACiht+SRcGYVE+i/qbEf8hAaHUEbAO1+WUv4kd1+wIU/d9OT
9KO+t1Hsx3U/WPsyGiCm3qKRKsb4tXRHDxkv5vEq4o14TH2JnE/nKpnradjje8K+5rfme9kbzEKx
Iz8/8tH8/TxslwDouJUiXyGWMC/xJkX0Fk7xmZDbXywip4O182sRtMlwmrJh6ExuUTkZEYyCdg4E
LYZY2vg0pAIoCJtTYI8OBQVqEplVSWbqFz1qRPlUNR8pNACeJzUD7IOENiWa73N+DeIRjKwKZve8
6Vtx6SJqs+4IhVXiIElotfL89Is4vjUUlFvoC/SnT4UpsmovlIFnIgAXPuZZCnyJVMzWsXG1h2Vn
u5uPpl+ISLp2/lp06bRTI1NHfwG6EyAxE0ZoqdQl9uOPCJ66C7ajyk5v+2uoeRqLfOJ6XDUCPQkZ
1JSb60URt/czR97ep+PN+jaCZbsR3QseF5RA86ex60eX7c4y/R7yb7mAxj8JzNYzjL6GuS67YxRF
UycSsf8eo7DmjNNV9gC/gE+txIFJ0JJ7CKJc7s3b+g50aOAeeq8AHQ8XaXzntcwt7pqvhWwWTvw4
5qKujHVhxBPKBHU7d0lR+VoQ+aLMmahh6i56oTEtU6TbiOiLIOOAiJ+g94290m6VE/tAJ4/K1sKF
VOamznJ66TmaIO4osh2CWdpgDrEYjmdmh1qGab0hMJ2PFusiSghV6OETTH0CiSTNJxrDjrrj/Rl6
R8v2/zuHm1G9d3yX8uNKIBDhjgmmEGnzFKA4d50/pjKcmkjDvGSJ5rD5WooSMPGJ3vW+BuQUGJT0
ogx/2GDoIWn2d/zSICP1G6njB5FWGQC+j66eqtSdkT++5jNWgAjCXukDY5/iT5iDoUNOyKnbSbyc
cMvmck+vu55orAimTQbvPMjpjwEzu4pOcBn3ejQafQQ/4WWg9c9TicSFJB2yDBlE1zAgqMLhmlAC
v5dxHkwixlia0bjNNjNbEPI+PemsackM2Q7arbkLeR4hgYCvkV+rQhED8MSm9ridBTbog67mlkKr
Q7zkF/NVSnTAGvFiSZU8+ymLSwCoakdP3a6El2j9yFjYqQq07N8/6Ex37zEIhXSwVkjADBY4dXgj
eP0Oq1egF5b0InSE0ldsoZkwLvVEqg5kX4w5HGJFKhSTM/tHc68RNLmeXRKHShg0sFG5ZigMCxhC
E1HfvAoIERkTLQai7DscvmaHmoqz4Cogy02BzVZ+Rqw+hiJIHHYreE/6cq0UOwrH/jWJOoPhXaY5
r199xBl+kOIF1Vdvr8771tOM07a4cPYlmadOHvzkbCRYfcdmL0dSicYdoisGhOSD+U85xSp+vvaG
K2zH2TIXikdWQcW0BwJzIxLAGVL75LLxJdMQ0cWCXHbn82Iw/c/Wp2N8VUDW75CcRrKTOLZBbLmd
o3lwlmD21RJBKiUTxl6MZtXV23mf2cNJTOVWTtIZNzyCI1k/IgOOwmbiK/36E3x4mLjIsY3pOebT
Yb0lFHkxHxhgffa1jv5eT99jAFYVq2sM/yMTRoxdgGuZ55w9Nfv/dzlCY9IhoOrmqFOLV8ucmUYt
mJLMHz088iEJFBkpL3HKpBIQ8bLuSx2w4uhYnTwaoJWcuFElKnjGtd64MCvScTfgjGdn1IMPfgXT
LM4G/ORmk1enffE4ISpl3lBxiYhM3NAU9gj4AlaiNhLi5fxAQ/iQ47NsWb8VA0zPQSP+aVDMp1f0
9KPvwu9z/lDxQ631MIiZSWaZR6zFNo/VU9be65y/7rh3k2Q1dB913eTcOHkai1LxvVuDYFSQjbto
mtUU/9gYjaeLZM2U4pgbP4rnfR6fwgQEap1U4/QSL1OQvVABE9j2YdOQ1ADZU6+LkAewRRWGnbFB
5D6a2PJAe505xV7AJxd3i4xeGfcJT7w602rrWOroPRLmFU5L35RqhTdgoCglbGA3vhv+kMywerPe
1Iejl43BUzna6wPJ0j1wyuqq6+rteHkSNqaAPI7rGVC7j1MbNp/3d5qEgMptV5hudnQ69N1kCanu
edAd0RTWDAhrum9hufwyWmKNBbkA6d7mHdCxmHExjSDi+MaqP8Y4aEU/ghclFJ57eO+2wFOfeQeF
8HKQLHmJZV1VpTQwrtXmEPwRUrWEkmco/P8M+YO8LAaJupd0BufCukfPb/LYjA9ct9UmWSVBdF7s
xR3iliCW+cgxqeOHYj2BAZmDnvwtiVoyDBAJzJytyrJvAtM6ZwAdIjWzzK9YGdY1BDT/ZyXW/WF/
oyHC3OVoQJw5knfxYXqQ516b1LKVoxzfeeuu733M/VCG9g7cqNKwsWIYOMNr/VIZFU11hppOIj7+
KCWbr3NrAPZ7PK3Vg7rZJVwL4ozygJm2DILo7ZTcirSLgOa4YGEJ8Fg3arDO/hPyWNIa8uTUu1u3
0dX/f+Pte0H3XjlGpRhWlEvBl3gYfdiVpzkox0QS6/KmWsbA5/F5S6l7bB7Yu99GJHK0YzLhDizK
DoTM9FyhXDrFRTAB2q4BLNjT6nz5DUgUIxrbK6EGeN8piPKwIaU9RV/Khjm03IJAYXtlewFIYgjz
KnGihLwNUeev9jrjNY6/ojEKFtH38fR+kn50qI4/puSdc3/8S17j99ZQo6ymVFRXSY/AfY7UuAuP
qJWg0G4EUEUihK6o97t68vDspjPJeeeWoWWvuu2tNpywlsFoKC31UvuC4IqeX5D9nhi/6Bpxtfzd
1AFKKbwWVfhvI/exDKvmDbx5fN4levu3qb3BTorcnS0qw7wzZ53dC8Pm3WHAC36iAEqIF7JSKH+R
k4niiykqj/tFM0OLP+Gh1FuKHgSgszH8j4J7lAukz5zCm+Ju2LaRh/hz3KEjypzYeEoexUUYH2s9
ANunDxlUoIhNo5nDDCCOG48BivwgF3Uvn63fFzdBSNZs4M2sQwbOpAi3FN5djs+30o+9BbzifhtO
1zlRhuUpkoyqxfEa3YEZKsCFUTb5rpHpmrXAwsGEC2sEK82wbBMUgCEfgkEUcHULMw0OrcFbLTw3
XW8fTvDO3ocRhnhPOWzjUyD/tYfthQ2/109hVcYuMOTJZdcPOVnjp2PfQk8aXWbSG3DyUruvSkFR
tFaWRiQwRs6hn9wdtUXZeSFmQQt26dO+6xOOoniWR5DEkocR3/MbJ7U6KWdSbFztAP2QwgRfCUui
AsBMph3PK6DaF78HnlJehvnDAOLvcScm/n3GbV95UKNa+bUjyrNV6FsS/mIw1WZrDmv7EfHrVB8D
A0iQevW3gF0pf1RgsqK7+COxoqGA+9aFz5R+e+f31J92t8M6793RKY5ZGEMVmRTn5GeZ/rvqbdxP
jb57aIfljPx70ATsmtpwEDcHWgpYIKsbyaR+lfixPvqh14JvySQJulvhfT4lvAQh7jLlLZXW0qjn
f2nYR2oIr7xMaj4jEg2INva4bDMj+4SPbL7xUfAZRCun6Vpmxt9miZtkahVEUCuqjFrEtCICC8CN
uTnPN2vj6ZfXoj42IAj6vtoMN0gqWObuah9rkJhRsNoAPgn5pKiqiAlIHo9Stwfylm0UpGYRAOeE
VfCkT0O2p9SMkaZx4SgDl/TWrDssycLo9UAOkl5Y8o+4KgMCqpadun1GME1qMVTGAx3YHjj3cRJD
PRmHezda/NvAq3OoYcVBPEibM9BSVt5PXpE9o4qnOZZ1NyzUL8mXti43LQPjaxWDeQTHpMGIbUpS
nhYbCOn5yWs5NJxSUWdnuMcieCe9Bm7s/7p9ydwpB8w2RkVO76VB5IDBN2RFSFscWOy5HNXsYaGp
gxGfKP2Jru9Xa0Fo5CzREdmliEHLLOE98P2ByooWBjAdMS26wBNReW7UAk/yzdPQ4VNRdhwXnP3a
mQePUU5Kp/zSKDyTuf5gmUE66jItitiQOQFd2wjNO81fxbrgQLVAOsgMmE/IfI9azZzYJoUR3ps3
xTJDWjrTQLgd53+6pYEStSVMi7cwErE8UTOCl4790F8G5WEYuSTCwPXPRwggxJjtYEdnv41MKTpO
QvMu3YKFexPm5/mCADPbHp85rb4KGQVJFY9haUU0kJTijplQgMTeEwrvl3sWLIFmpkNemgSkGTh7
ui0OJARPupd574tFfcTBlcgwVxi+2Sj4ipECj6ezsBtcwCzm+dXgXWHoLhPbiQZZ+r8XhnVCaopP
8PNu+QVo5lK5xPkPsVzSZ5KcqsmBO875wMRzRXrw35OhMUST0frE038gaqbIqgMafzQ7Z1uhr7Nj
JHCAgDFTWz9ibxvbhLuU677EQeU2EmQaGN7swslQkWpBSj1hIGZb7CAmTZ2c0DyVOq1bfjYbxD8o
88NpprTN6ztH3Hm1LRKUMM7BBBE9Ufern1Es2JntKHukHDGMqgYiSCcjkf8XEQX51M9V8GCEDd7b
P88eJ55/ev7splHs1+CTML35V6IqEAvGXEjLwalFl4+FsarIu/l6AyrRp2rp0kwEGrmlHN74bv1Z
/lRCt+rUMDsjf+boa5Ma7B7g4XdzInmvhseuyxMerPvROoYgHvfkhHsvPU62rEhvn7cjjXRkfFlO
ssI6vljn1hfc8GbJEajfmSjjCUaKIVPV9VRlcw5o9cMhs0mKYy6QmiIB++jFbdvut+NQzgL8am2N
BuCR8fejHmXiSsw6Xa4T9G+sK2tMmOzhNjzCkiTgitDNclFWFBuZYoUirxGhX3VHT5UfPxy9xbj0
ocK6Tt95qaP2k2SlVKYWX4tSiQZJtdi1bAUiTY6cfb6Hwa768PbdwYb+nZXnL5t5WdFhhhMcZK9k
wKMNzu319apppdJ8/9Ol5Fz7cxwwtQdgB/XY4Ta/mI3J/j1/Mc12j3cEMG2FAq5fFxmLHVDt4oXn
zlIdnG1I0u4kwbvrB8iKXxCy4K3NO2K9nSHV5LIfm0+s4r3TcydmonjUmvu3/pFYqZCByCLoDnvZ
L07+ylmGWQK+DK6qi7ahmqypurvpYb60rqhe4GB7KlltQqdc5+5fUvp+t7R8vFqDhl4E4apeG0vc
UoSIWIoI7KeGnpPleV4DHdq7uYy0mB9ZtONcD5lgpETJWYIKK0FfMwacxEJqKDdBL7qwzdx/l2Xv
R7/s1kRVaCSAqvlqYno9mppLGhGm6DzzSjGrEeIZ230NfYPed0Dipj+1lbYkVDP5xlRChpYQk2Zi
GfDusKjcvKAP5GWmGBe+I4F021vcdcvXhSlptPXEuU0he4VyHZ/zsvgugTHTQ2Axz84saWcPxnzF
DilZV5IytwJJzcmQ0Q91ugA0X19VnGPNtzuU/o/WCXDRO8sI6aU7Onj+xm5iK7Ct+Yo6UyyXQ4jy
UfvbWwhW4Cd6WpCMfHHtiKdizXklOLZ6fvy7Jm+omxfv8fVmFCSCerbs09byhes8IZTPvAK147Wc
F2AXZSUe9aYAXyrlzdQi8avIVeWZmaXw8yt+cAh0lnjjZPaqxA8N2x/IzvR/C3gg1fHT4OiHXRI1
dXOVgoSb8U1f3lLe3g74DS5ykArOQjavfl9vHhOmJPk4ggkpNIQV6Poh21CEsIWHHuDzWlcTNt6C
9nZ3ORJV4lwHhtnKWr8VPiAg28sleRDLqMgdEoUaNM3SWV5TWjKh3A7zujWaS5uS+72LlsW2jxHB
8tsy+6WDlN00gJReBM+ey3Cwe8KgpHTKJMugw9XohLnUIP2N8qTm0nmKUBbUB/mZb/Mu+lGrPz6L
lzQfOHilq2QIMZw2JMoZJmRZIw7nUl+d4Vdnw2exJVObDzdGPx8RJ13Wj1QZnSck5cuFAq+yjv7p
qbpQ0Yiwljz+Ni/6vYqorrHn6Q0RoEfiiebjFHFr/joB5t5OlAgahUsnwdxw87ES71btGCd9Nbwy
z7p0qedephBuLRGTdkQYSldsEtufMmKdOFHNQfK6CsGUHB3RPFhv7KAKPXA2SRELoEHS5W48W73n
T0f2El1FjGnlKlYVHXbgpWnNk+lyEXKS2mYSirIjay5XMx529WAT8bbPupxF4VostaWbnPDefPvd
T7+rzd2Lb/GoR2kmw+K+Ua+u4soLic/uI+0dGGgomf6vRfHY8tEAYZ0k3KnvaLIVYMlbmSYD3t8F
suqB7OvTJVVBuyfnofS4fgWRmj7X2rviWkTvs1KpiFXFcCl/zpepXDDWgy5QfKsDux2w1JDzVYqb
Q2iVUei0JaDQcfyVWXtuUpDMJ6QN/dl1HW4P1GHhsnsBKC+WlL5dRSJNxEKPF5GfLnatzsYG/a5R
KmguGlfhrE8LTtsUYROp1fJxbtCSefJ7wT0hdfwPTNNnkgWVdH5RbZY1d+DLIkIYnC2tXnzllowO
39MU0duWP2MU7bRHQLVo6jP6kvQUrOJGAhSlkIfutzfbd5vAY5R91+H3WMkAZDIRDT/PcBVZevmE
jqVkMBjCAl9f6Wb4JmcBslc8DbP/4qHd5olNKckWnFnwWjKFD6qph4a0VUeJJ96mbxeNfnS8+LWV
a4iJa2ND8M8HAEcAlrXBWYEkMblQs735HZecM/gQWfbOZjpBOcJqRFC2LK8v0UogPqnFR8eyMEFc
QDn7yX6gswEVTwI0i8WxyH8Gf21BTXm9my2PUhArXQr5SN43Et6wM0y/fW/qx6mGmPYatq1NiSso
5Ekr2MBt1p2sViTVNeW00/r4d8sDbiolc34cKp3bVQfkoT/tG3YSm8fv8DFRqHzxDC7k9oPIez8/
bC/EKYjBGH/EubsBmf2+aPKpBNiBemCHVc93sjOJ1vpNo7OI00MyIJCrXBP5ci1pr+dX0j6+MW5j
pWiaW77ErgHELerTVXBkwg9JXykmhPv1NtMUMujWmpz6wtSWjGnfF8b3cSCJE6WHpSnP+7y7i/fi
aOZalr1dlN9PkeAVc5JHWi2jm7yeKotN+fTGyMXjzrTqwGFhwXcXZoW3qT2PWaf5mepi4BUNPjng
xvDHFTi7QdxKJ30sgk/ZQKmKYvDrAafmBHdd6eF3IDS/iWVwiQQCz07R9o1V8PR45Mv8Y2KM3NHl
DkezmGYeMQDlkO2gQluOQwru3ZQh429fZoXl/iDiZHIILJVEI5U6sOCn/O+i2UQPJhWKZMPuZYna
E42eun/3tvSH2v1qhCNiJ3hhdUwFLCT0hgXAE5Y03x4bviqpZrCzgufvro9P4Dc1cENIFAD+m7ws
kmFUOpwcf5ktLWwaOa9ZpaAo8mYzppeRz+pbgADJRheUPN+KcJ9p1x/PqQvE1qvnIunJm1OsZuM9
qEF37FtbOsOdNyRErn1wV2uuakRC76551ewtFczRpzH1eCSH7JAd+9Wkddq8nXVlMfXsfC2C9zXr
Nrer43m6GYajIKbHORzZOPFUZsGpjGgSJDzuLGJZjX3qrVMqKFH+Q41k5TgubO12rz8zYd1yIFve
VcFh0HIOigE5e/Yl7+EIygHa43TgDugRP0uLBBjGhVZrWiePtFkO7OJmAkNL6hRRKMybueSr0j2w
mzzyuKGi2zc8uNZlGkjgQXavjWm/2I5VeSobGJN3/TXCsvyMw67Dc5AuW5OkwJ0LXLVjcv0KVHn7
2UW2JYJ4nkUXj2xanNmQArcHRMsqmtI+MfLWY7Umz+aR24DFQyljZzUkHzJhjjitv1jeM60lym3t
UfqR/2ECBpOTr7gnbohLWVRPmn/FJgBwVKiNvv+CaJOOvl8hCBU6LsQIuyJDExRfwEMQJPf/lJNd
27AXEmxRLJ4XH01S2wkQ5tAIGNwneifD7hVnUC33w1k/TQf2JtdplJfKooIayQSC4tjyaI6gtK/J
ORS7ksxqF9GnSdNiIbG8FunpCTlrOtqekqcEE22Pg/unNYEyYQW+pDamjj9gv/G9sx/pQLb4TP9I
yLa0dekySRnyOy/GebBxH8r1/h1SPZspnE18/36iMDdokMWy+6iwyOXjlG44C/0GxSEizefbE3bL
ic6bUpNGUOaxU84O/v6RjUZgIQSnZGeTz9idKK7/AjNP1sezE0IELfIKaakGgjumOmloRpccNReR
kN2Q+r5NkFrCr5RyWl8Jzlhs11fvx7D+UdGq5KslQMk4DvJO+B6rkfdYUdPH4DCmsYSC5YmpyPbS
P+PijXd3ERK/H+a0CYssTZ+j5+8bTiT3n7BwPAETciCm6Pst34orEyEnKy8+HsmMNptUFfkZITw+
7NsGL57GQQoZ0tydA3veFrOm6DZddlBF6Xdv2kLVNI1IBPKdlHQlqhKHb+3J+Qkwe0lzBbXEZ4dN
mcuybCANNenEN5wPHyEMf5xZ5GefxMMRqqQtVuVnQwxGpohgU1vfFk5CJKSvYBxxX0AHJqcS/AIK
XcZje7u1zp9C+5tmSFow3GV564eO61NqV75j0QDDob3MaPJxzIZ3NVBTj86wtMWA/rJJiw/i5VmY
WMr2VagCGDMVqGaGYRf9SFJ+AJyffjpLn5XUqQE+s0QfbtlUNzqZZOex4rjmz18p2nZ8yQiTCh+l
Ku6wRpIxJkOF8RvvVsnIy/CnMHMrUtrzgPA0RLKfz9YuY29qM1USGaNE09+f+5cES403PQm7C5Tq
/S7ZBiA0OPy4SBnKAbSV7RcMXlRlo8A7Emtguysf1ASff9NlWBLm4AitruChuTju4FpOfQSbOAjg
PjCswRS7K7HvIvLNMCBeOoddU2MTtTnkK21VTQdKigL/UqYgqNWoiAeDNh0Ku6XxsUpnsjCH2cjW
PdN6pvsW6dxsrlk5tWEsv+AYxArpuQUaHfVlcg8MCGrQf4x2aRyLP+/Etk1+lboq2LHeIeykX/rw
m+8/jm0vLc0r6s3nY34HUmRlpX5ior/nIv2oe2gkQM1t90n6kW8TFpO8kJ8gGyfumTipOxf64xCt
5x3LvjvwckgxF6YcsriLT33FnlG/W07t/iLTLSgjQTI/22UOR4nExyNTGGlYNsitb0UhkVqE93R9
QiDfJYluYJLH/sogb59jDe1Ipeqs0lwqI98ttGLc3X0FDsfnqQWdaYp7aSzpUSO5IHp8F607YSc4
TbwYglR4o3YViawU/Jv0SAL1cCGGuZU7yeD/j7ERKal6lenjkxhBeBqVANcLY6VHiuEB+YIPABR7
fTPnyIjk4aZdvwUSfacoHobGaE+hBFjErne+PEOkuHuXzpK3w3aYNy9JiYfriAn9Y3UXycJMdp/X
cVbQZ76TSa34NIVtuHxgs1pv4ynT8Rkh/94sujEN61th+wufBW1srhZe19UIWXfRr1T2tYT3dAok
cgC47abJnnOfrsrkO95RGCOVwnSUzbZfthS6qx761M2/Zfpak3GUx7lBWzev8os8zTNLGS6lqwwT
P87ALWVRkoJD8vYuwiXtdqgT4vJUfmnB4L82jiBdnJAKPDMQhDwJGwCjbbm6kNwGQK2YeOkaMsFx
4tkqP/w402UhRqbLILf8enEYCMq1gh+HUr0vF0+vTVsSEzPPlnZgzrrWzrvO0wqOcNpntcIXKB1+
3G0MVEeApB3Oo4KuXOArlZbWX7AKXmRCv8Xc2erM0TYnKUNr4IcMgJJVY/argDeeFIOkkB1A9kFE
YWSQ0G36EUbJhJuDusIXYo6rCkMuq4BhMebteERoScmgk0zzVxrK3bHfgwZ5wvBPDSzxQgcEEQhX
Byf8TrQSppLAeQQ7Ln5kLDAJa2PeGcZiEZfFWj3sFiuv2BiB2snj6v2ZSVWq1e7fsqGaoXPF2DND
xMliFwtSKuNA4qhmBY9Mrhlg5+2dS97LdEY1zfXqL5/VSfplLSiqowWydUadCsw5wna38Id4emR/
OiMkIYysUjYk1baZjuAgmZ8dPjBqeSk4OVv9IRjDcLPVt5HkA7BNsYr4roQXRXPR4exhBiG13dS2
Y9tSfMYxntnc5gC9LuZqCkVDSZgTCMwa+d3YKPVgtFcDp0Dn7BE3MqTDxn2xhwNBx695OVvnsVu0
6YynkeOWJTze7PWG+nOOUD+dGeAqjsqVttbiLEcP5GI+3GcE14pgP1YqTyRT+ylWMKz587ZYAyE3
lBlFF3IUdVBRthyzrxMZmLZtWK1xYpWTG1W0YpiR/4AgzrNyfVnZqNTm5bpaKiHr+OvChY6c611h
3sCBvrDcf3nbjEiNdNz+Qr/r3OBztgkGlrCmA5eGfzcF8EVUOZRs/yQ3sixnEu9YKm1E83qV0VAC
0dGrVpvjTXCDhUjWsraGuDrlRWDs0nxOIcm3EP2Xov/CBon9iQ+hdWDqgVF9wu9IjA5bWLMhemp1
RwG4qeYMeDn1SiMr0pf9QXEJsdabEBXFbkvS7oOjkqAqbg5DbiWQ3JYf7wJN2r33CRkyVzvHTRTG
hr1u+7IhNf0fMjF/UDLlT/g15pXLnL3YwdDSEDq4LeJfeqgAMKJ6R9XvExPSjzEYeAJcfyVN4XKd
ZrZdLYtyMMBgn2QJ0/jKw376ST6aLP/zFkTTULpwgyVchZNJr0L9fhtZBxohj17LoS1v8o9QsGkO
pPjz9UanMA7SvXhOtkEBTvbKLMFnosnvEXe6CjySdDecs2uDtcylCYSpOCTPeYqHFFxmqydaiOAR
R965ukyW9f/AB3zjhKBdz3hwwCIiLJvlIvVW7sSI6owmztgNSh+cEzCw/MpjzYaQt8ExG+z1oXcS
qYsvGYb0SCPi1Uy0I2VAxF0CBbh7rDXea10p8rqCQj9CNMY1N5rACOKOmli+GHzCQWSuKpmD4xvE
9+7TfEySsGcwUpbikMkMdAwchihAhI0kafQcU1MFiHzJbFKpl9CC8eiCcJmzUQTK6zda1S0EFO4u
a1CV2Ky2nLnCTmTVJipu8d09xfvh44HeevpfZRklWEME6bm6aAfgmIPWXk2lFNDAj3K8mLTW80kq
Wi9Vh4nHmjnpZ31TE2d5uwO2+Wh1gFMTeSs4yIVPKKMXST4M/TvHeWwwEOVJ+SRbVwh5gpA6apdx
Tsl1EHls0iUOZbyp+zZgDeNT2rY9wca4kfmXfwh9BobOBDDOHT/uscXJsR2pJnQKXqB8kgdBpJGL
Wivq/Wl2auWoPvA8QEok5eoIjWtY63Nbx/TAcFPCbCIxAJVKR9gwAFvpuZCYErUSjKjtLjTmHvKp
zOkqOVAgYOXfYK0jZf9EYVab+knzHbUs/yBC53STK2LChGoavWRVuxxaT09BYcRcr8f+zAvyZFnC
P25wnV3uRbD9jOWf69Cj+SJNGstH84cqSVIuklS/6G97OP1aY/uiRPVRYdWae5jmZuZmdYsEKMlf
ZUN14pbNXyAssF2fANloWl8Lu8+DdCmbZhFq71mVDypOU2G/B9K3MjfRJqQnW5nLvKdYaWkxbxYK
02lpVmSqZx+Y+3i6rcELC0R7lo7DPuWC2jVCsfkggJ8cMg4HBxkgWEX9Mo1DsjL71BRZ0CrdBfB5
2pBT7nnAp2R/NSZxY9n6rlS4sBu814n639qTuavvd8TAZqw4nzfMZQTk4jL8eGLxlB8Z7Wvbos1u
ypj/Y5NeT5ZSRawTX4Yh5X0x51+dlSpDqLsTmgRyPg7vaiyG9++aqwEWh8rIQoUkJo3qyHH8A9Jf
S3cvzqj5Ditcah9FVjzWhzY08k2thUSyWpoqUA+WgNlAzbV5hlyoygiM/cLUGuYJ1+GFkuq33ChD
cLwrTA/6SJR2r6rh4BfXaBUHdW7Ze0oih5qS7CQl/0tCqLQODdzgrcigO/4aGGde4fZ7tJbt/4ve
TVXNl4Ci3SCZ6/41/9TNnBJ9vquOeopBONEhADiIJubnHtGgLNqTFXc5hNuuGxMv2yd0UvjBa8OW
JxhOzSoGAb7fPqM3iTLeZZSPIYstGKdxAA803kXvcHdgkafkgookvQAjU6fxfv1NdqwmBg+ggoxD
Vejiant87sK7Nk0ZJzNOQMojc4nYXfMX4S6qST7NSKiDjxF/YQNWC1EDjzkVp3OER9JBHrXVuOpx
Pu8dwsMZcScG4GtYlWdIO1UE05HT2HtJkP0ka1WH+YpNNbES7qjjNP2mc6iH+j/AXf9hKHP6jS8N
YAv4fWPMgRdNjGb/TUn0FejxzlDVKtL5hWkCOPmC+G0tf8cqrg1PdnMGt6PGpD/vAIT5/ezPdsQe
7QD9gEObAAXIdWhuf1+0A53cmC6cH8Hm5dgnw2RPX71FmTEtrdutWcM5JY8l4RPNwotqUsizCbMD
rF5xis1n7/V8DeeS6R1L4OOjNnYzN8yB31n1tOWYcc6gowzFop8F8TxJz1WN2A+IXjkVLzaLGCI3
DebGIwx3eXge9+OOyKiRdaSLdcXLeVpv0GdO+andNHstrhhfgKSDzxcK1/hv64s+gP6JE5iQpN9D
EVqAdY3figQzpYVfejRAYEJgaXhW3+wmTaNN5SLAW4iESSOuyTO97zMdtkva9r3C+0r9SdQF1buy
Jn1TRBYdNL1kprIoqySHzmdS7owwFsD9HprNA4PZ6mqmE8TezkJm4LIykYW4T92nFO8wfGnyWvF6
LZsLM2jq0u81CL06Ky2+6ZDQFdBIKg9tnMR2PF0HGfoR/0TqHGuviSqIl7Uq6gS9W43y8D0pkWmr
rTg3BqjHxfCRbtABhqVuyFk/JEI7ugv1UsrZqz4XFIyUvKooV99XluzosSS6icmvdw6fuWRwLlrr
dkOVtUfNSnWJ28INKWOjyDAS5u+tFWutE2nDiItaPP6/bvm1fZSYlBGGGwylbEEwpPfh3ISV+LSv
AWZl4C3Nh8aq3aVOPdn+/ztStFGVJMbVTTyrrkr9g+zuP7cFy3Uz/YBX0iOEgpwpx6fUt2ZTiuky
ftu8fyKQCSJ3A7NBMWDEiJPyH1g06AhQVLI2+90klnjJkT9xcI3Yj7ywz9GS/6DweQQauHBgsYRk
dcxbopstCqdRyUPsNbOJ34U/3tU+ZnuiH9/Es+vgN7ipaab5AHIt6OtNfIcB7ChhPd3OosXQqRKZ
2D5AHuQ1w+ezlb55a8BjveC3a0HoDID66fgegSeBLZnhiVvcki/gNbDIjs5RkJ8o3/OkRQjpJW2Z
M91VOCXX68EbNkts6MhYWRLM1b4a2md8y/mVJ9LnoMtVeOJhCCZXDRduCX6SuGMAG8ma007Cvu8J
Bu5SgZRL5N581fx0wXvAofvx47U4NWuZGcW+G+LlpLhRxiqNgpB82SpecTcs+L753zCpuGRwVdWo
GMVffNMZC0xR3HCFfKdNp1Q66sSz/UMrmEJ2R0uI1C8db1+YhXsXV5xL1qUZ12TZZDs10gyTHdgJ
GhcvxT5t2wZleEoOl25N1Zt52EYsM2UVBV341PBrRQ0As1tpXY3F79QUzzX3HsbOD8oXqyoiiWX6
KvqRHikwB4FpedlKQfpOwn20esCGTxEmmgTqdGCK+RlDqGiYt4JXeB39piPAkj1CTWZz56fGDX/B
Yyp8mt3Vtd7tZuc1VGkfBZ1NxJU42phzWSLYQNhS/Tn0KVrYU7Ya5kdscgqK16KPqKa/9oD+eL+V
Du0SOnpBQWIq/zUnXITvbr4vFJMga52bYwllpo9fNXwjeJ5+0VDnF/gUbTILuFocbYD3yyH1Mwfl
ENjFNDIKkXEZ+RO1u3hIl+My+poh8YUg0tK0PlIfLaafPzS/LrhPNs621dMQZ77Bwv/bel+vpFGH
WCN6zD/oEBTBYG1UL/f2ppEPvrD2LYkN5fTBomJS1gB+I/w2HuWeXP6VxKkSyeQRUvXkh/wQRQH1
nWkl1DKjj5BWDxwFLbYX/IkVQaKM4CdyC+9YG0h7HPnswkmhH8HUVbuY9pGT3TBq6kU7aGaivi9f
tnjuqBRvGFKABtn8mVO50WQvb3+rT66IUEeh8hyjiffGaHsdJ/FaHaU289HJCygjejy1bbbeMtmZ
+g20l0kX6H+nuVAHXteqAob0CYXLJyr2Y/ijfEFAfsviKSwP7VCyPKRzGKWMHtbToBb68guWBEsM
YaqD5dvKZ3TZ+Olhggn3z34u8BOPEIVdTOhsABbQTfXeMlSwhYUAfQlx7k2W1eehMg8SS6LvGu/5
4BcmE/uzYLHmeGKdgT3V2hdLM9gYQtIqS8J3A8Ou6vq1zvRsZaCk/o1lpznJqmkpB02eBk3i1sZu
MnjLn0FklBW5db/G24kduodMHAcBnCGBMYp6al2NvFErLc7qdoheXLDvotz5pCDRrBDU0aOi9ze4
UlqUb7SSEU5fRLo+Tuel7ALkhDFJHrG8CBWc4YRograp9UHI4MEjNsAP9zCnRfyTZCDQICFIXhUS
u5AzqGcpnMXOL2En54XXxqCCs8DcWu6Ka9bW/1kiVwekd/KuJtkMMf6w1h6VuuxFCQRCXj0974/V
OiIgyrRWpyhT09SyHjK/4zo0l6bDwIuIJmq0TAaH6zJMdpFHtSFKGnjR2RNBA9JsejOaRb7s/WZM
w4PnCrrTvXMcDF919kwzfl5twYtLcikwY+YpmTsuYSocFAVhwP1+AI+tR0+eHkEywzpMJ9RjWH4L
clhot5UvnttorK41tr6aGwEZzShvyjTDBjLeKxCTn6t2mvqaSHNqQ9TzgH1SM6ylUAjDJSavP/dy
qiztYsutpIE6zi4Gndck2NjvSJCQ3HBNsmJt8KKihSiNv8G+FPoN0OEgkPCfwgC2NHwDQc5l0OB4
aT+z+5HJA2Azs8rf6FXKCF5n2K478wpFrW3KTm+g086MVLSUK+Bc54UPFmqkobfnVIVwaI2LdEKW
dez/b1UeHhX/NHGECP6cHmqCjl4mcVr9jv6SSkfGOo4ICv4ZhVqShChkb9dFslIXVv0dZeKDaGJx
gxakLR8a4QqN/2u6ZzgFq+6VpsIaUpQrdvhAP0dKcKhyT4Y2DDumS2nDLMxjhapTJjniVaxyKvDX
49VZ5RKykr2WL0TNx6T6bVB1FvhGkJ1Ixt6iRxIHnI8yoQE0ZwVl2hN2SGQENge3dWGTOTlTe1gR
3B6HWMDmfR+xD+BUyHjMhBL7B0XiwgagR8Nm1GSYH+Zj3iV8JAhMVjYhL5Fxj18QUAm518mLhxnt
HPke/Ay3XVAx2CJUzCxBYdWTbkKlbocURWYk1gKZ5/NpQ4fmzDQEHDUkFuYydmCMLwkR0e2hKZW8
vTQfM5Mff1yJmlto3xxiQt7TQU0iVsJk8pLGIprgA/xbL+MXjo6opAxeXMZIjecLUMoVC71rMkgw
5N4I9UrLwO2lMHMal+hc7qpsaiTuXwIJZxvfWv8+m+s/aoPgHBrNlKpH2ZMqOc/L7l9snCAHb9Jz
nLI3qnOBDyJceeXMBbCpHIHTrJJE3aLf7M8zwcltWZ1aURbn0i/xPXZQRCi0L8wpKwzOBeQip9CM
Wx1HzVvO2fw3rIbJk719QOOOY3TIB3RUrYuciD2GOD08pTkMrJ+fBE780U3WnfayadVCLbP/Wnss
xdxM63YlLtXWlj05coCs75Ce15wCOzMCqt3Zu+JpHMM2t5QL4VtETKV1lHlTbx2bz0f9cEvN/ZJo
LSEdQGRLGJ2hXQt20MnB9WDlIPDC0BgM07mZRBx0PP8DNonvsOfDtpgGUpvEtv8LVesdUJ/UwoLG
hUdYj+dPsDIpVFHvQmgaZkrNPDS4+LsOkraZJ1quP92mUrMo5m+OpRLVqBVJxwcFFog/4YdR2o9I
jBKHjS+eMVcxfAG1ml95n/tQyKWADgZNgQCxIkL78OJ0OjD51EOoixA4jLkT3yWYliwg/89yEe+F
6Ag6miqUgqFpLzqfnk2Im2/xIxhfYI9L5lDy5cP1pWMaBgyWeO8CuzWVwuZEVXJS53b2nKL8n+Dn
cQcEwqCMaHyDc8vPqqKmXqBx3woP2dXO2pao8zgHNY7XNEH1dTJJYAEHR/Fd/H6lTclhusGwDjQF
gUEh4UiQdb/nGSBZh9pzLmPOQqXF/lvLFW6SUu4qqr+/lvP85CXz2xlND9Y3Zq0ckNMjTQLFqALf
0PNg7MPzKPddDno+l1qi9p2lqZkaaJE7TdzGrCmdHHeGaMG4kXEO1jLO9TCEe+yJi1lmExIJsiU3
ZhN7/eKBjp9a81bFm15LmurQwARol0DpTWYT498BnXD9nhkHjl/mpF6mNdE75nrnXv49Tr5Zeram
fut2r1fJTcqV2Z8dRgDfokcVd+kQlUxF9bTYGbVseI/Ia0aEJSl3v4zfcCGU/yFd8htGfJecbzfG
Tgxv7tkQbsEwMPh9nZ6EEK69j3Gt6qT3RLaEszCapNFoismoIF8cmPv4VQN961izFSiFmiN7sOFX
80jqxvN49gYWo3S1SWNfMXIfiByuzaK6YTbj+Du5m5O8mGz+VXf02sfDs77t/TUEALzLspZA8Zlf
DFdaA77ZUjmwCzahIi4mmuTU2YF0hUOfucXAuBxeTzewb6NXku4aGHeg7GxrdCKxOxUeaLiTOio+
CCYzjn2HVPyrN6eqt9GoPB9AdRYHoC5OA4fS6FIAzjJMGG0pO3ASYhg42AghG3UPOfGRsG5kxcuT
LVAO+43zezGfGCKDJA4PZ2N+RVO6U4du0oUTufF0cHTbGPlIhRSCIBMmbmMHQyPZ0dE4lmSCumPJ
/32MhW1p+tkiZ8R/HVsm7q4x7wDNRnAm7/N3/2qb03vJ4o2Tj906ZoIxmWMMHKC6UY9kWXuRd4vK
ADPxkXORePWjk8Rnn1IPcjyRrVerqlFzFsUKuuKFTUNU82sohaUt7F5SIhiARUxmGKT+IuI2+tj7
kNXzKD7xqiMiDij2pzFef8S5qZRsZQ/nf57l3dk52eBXbF6I4Ww2BWR3m2EatVZ7zLA7IEOEtd/S
CRhvvgWK39g1uJoZDV0ydEtPnMe9GvxnBqwHNaUtFKHj2aRiyuL99+HCh4FOOgEdewsYHWwU9Y3S
ItOnYl1E7GDMWXDm9UeAHe5ty5cT2H/X/Stk7ga7lq93VxeycDkGJ5LWjepdcKlZgZtSoHXUpF+i
sMk9TJaFsVEwG8DToyk5nqSDEsaTWj7VFgSdS6eC86r/uYyEBvhYnTSu47ViyJl/fxte2WghcP9Z
F4nOYiKYN23t8OPYwZ4bNrnh9Na0CKHQAikFGef782Y2Y6z4xtSN6RrnLTf7sDyZLySo5FZVrqpw
vEtHZALG5/w6NKLzFxYeyJzUXJcT6O8I5KdgtR1tQc1pRDjvdjOfzTbrcCYeFuBaQ3EqTpFYUWlb
Op50Dynga/R5PMcVJZqC0SKBmr/Rm9VMt/3Bd53h7dyDIm/EQdmYqtFWovD7PjomjBuE/QPSsG9w
GrUPzPDR8SIvuulb6xZjWnk+2LYzaY8fmpfj40fLpg3MhqOoY9Gy06nbReyWTPncJzg2LnLvqk5R
IZuUksJMvHGzkSmQZ/hX0gES73uMcyTi9GmXoTt983PNq9EaVQ1Nvl9JeGMaNdDjWIj+rm6d4UcK
b9ZFnwcLZx/7reAkeWAlR/1jLkUnT5U12PdcdVHwf+q6KSinXFJ/MTB8qEeJio8kviys1vf5ESlW
Hy7HXctVXrg3mWPkMnAypE0oDDOqrSR8rS9/U64NSt/O99UsBHrJRq0AR3nb/VrYqGLjxMEhSdws
nW04p+qRkCpfK6Oz1y2Bhk1jSebD0Qd5zUF3CQpFVRn4i/01Gd28sOCGmWL/OBIVW4X+Faaez05t
QqY/Id87aujVtfSvYN6hBFPb2479UVAFi7+6s6tDgC8py5NjRcIiacwDZFi6Jbvs0dJwXTs1Nv+D
N7Zo+JQApZhhuQBa72rGakh7W83rSFWcefzVhkoGZWsYp8xaaE/2kzioYTkcvMYzMRfTr6XqVcGC
+hGBdW+78vTkKa6BgOxbfDBXripVjvpKVJ0LBVKeXTsxVS9g9qyzIYg8BMTmX3jcCiVgyipy1aIj
fTW5sinZKi3sPDWFe3To5axNAa03X9bpxoZqhlEojDThj/5aI4KZ6u/uIrR+OUPApVih9o4G96Xj
SePuVimH68n6zSAoabRR4+frsDOlych5vC+UsPCx6V3p3RwpYl81xrOOCh6bW9bFPHIMxzo6zp3o
1aTx/WNxwW3fR87FwmWoZvQBE4Cx60ls2Y9GvKTrWsT4GtG+hSsAljRUKLJupUppmwvQrrTfs+6V
LNNVqzwyQffuN4hHU2EX2Vcsr10pIqLsXSqjopBQO32+85oiTlMwP7TYSQpazq6u9X0DwIBPHB1d
plWyzonj0xQFxGcw5Hhv+hb9bgEKsTHxOkLcPrk7zL9oofGicP/IHuoiuX4eDoWLRM8310uctuoP
IdYiGde4nEACx+GYYGdH9Cp0WtgJVpXXuHs1/S/7cHP8BqpNDuF+HSbBczToRQahquN3/EeXI/DI
/MNjZBolEX4NbqA/c9fxjjhRdvh4SO5O0b9/yoaeDDWBbpjnIXuPTiDsYhAkfIG+QSooGI53sSzT
WqflF8OczsZ0Vk7F4RvAGMI5lOv1epzc379xcoRVbJXZHew7EH85YRNwLDZieYIqXdSCQicLeY5T
tUYQ96r17d5YeFAJq63AvfwHQr4lJSL/q0mVQOvBEvNZUa2p6zCZtqkVgVfDkyKGUFi9ZaUsBxt/
OSsOQdtWzKL1WCXundIzkwEL95EDGYx57Flg8D7cXVxOu+naNsRvPeeSHQlgreLgGUycxS51Izgi
CmOMpR6CMop2GplSqMH6opw1OTNYht6XRqlQyLoHj2z2RJ0KfYpFRd/2V2C6t1zGYTYwqdl/gCso
a/Ko6uaXdZA/fr3lnrXNP7CSNPbLHTrCGIO/5X2XI7zx3YgStKqaQAYBLfQqVmiKD7tmm3l5SM/p
2Jk0mAOor5WCcdHBagaWvGLOYgG6HwiTURXBPMrNyXz+b1Kjajard+MQ7JVc46GnjJYCTk3X1RFf
I57QDEBP0Jy71YHXJfqImmXufCQDCO80lEBF9L5EUAG1pAk4um/tzi3iWDYfoO2Dnf61LZKqIJCJ
9YkRnzVG8UMnZYt5D9V5TOJEeJEbH/bXSDOpuWU32RlPyhF34kioYjgb319+LTRfLmX+NX6Y97Al
i2uI+85zG0wMX3+BdEqrC1kxx0ZUOmExS13frL7JcrFNm+qMIeeVsDGGTe5T6YdaQHGerhaInBT3
GRfAWoE+NjoYYCNuEsXp0q0D8c9c3JzIZr9mPUH6xuxZmoRenaj7tjvYKYYCqcUl3hVQWE7hUg+a
++bHd3KzA+Z7IaN8HoGUiehCeveTmITdbCFZ+NibaMchJIwuWf2BVbEOb2AW2AKY0Qxc80sWUUzb
MUyfoEf0iCLx4d1HumcFwkXeS/pE5/Rk9mXs9Smdzk+P61xXQ5M/hLjsRFVcj5CPLXp9gq42kxVw
H/YBSnfhd9xw6Y7O6UUG20owGNlPCHnsvFqa8pB9gcykVyOwGSmmSXoLzaaODCeedjkTkA116Kk4
yExhJTOo1bGZ4ZGO4HNl98l8wRDgf3NHu3QF+INLDEjcHxXVMBxX+b0uLb5R5mC3M/dbeYB94lup
q/YABZGIX4Jl1XIU7wtlqqOa7pu5lk4f7hz0XNUWS+4Mo81PkrGskhCz8ToLwlNf+fOXwj5jZIIf
10ID9HS3pW892kTSrPFspOQYQaiLNF/IQVgGWkdUYSuhmNv/BHaUkKOT55X7Bk4/FPPtrL05LwQP
OcJfwxxv0F4dwHYj1ZyZbjhGo8Hfeq3eY/3aKLVKS30UDX5kLktWKTQ6IPSbmwDcskpEkLSrgOb8
AeJ/TVj3gOatoiu7B5DVsmfag7i/4jQbxoB00O1JwUqqxcrLbz13H5HcgsRVEAHIlKWxL+HvKKee
uJ+u2SJAwG8c0JVSzW0eAV88u7gkQYvkF1tofQRLoOS5tevNvgfjsyeIQFZpsfJeF56Zn1evn7vZ
05unuq3Xgt84RU9m6pV9WgJgaFN+/vYu5u4OI2Q2Nz49nYVhaEtahnA5zId5WOY7YEktXI20hazx
TbRJT4C/OmahUNOWVenGXJe8fu0hBi0IjruwuuOabKNBwWotT+s8guxgeBu8UPqFsgIUqjj5138C
Ub/W/7tjIfCQ9IDYimhxTdCb+t0g5ZOgDVIG5tCBQoyvm1ezT/dHWnl8JPNmqGxm3FOzEw8rGgCl
lBvk7b4dyadp9XCtQB35QICLvo1TFBaKlEgy7UdbzbQjJ9bOPvG8gLqfakllO7+Xafvl4XKVjXOc
Dl11BantUhnnvRYEiwcoyG5ZZAwptcza85MF2/rjqOcKC4T6a60yPJ+irtIu5VQHxtEy3AXw3hnv
tD7yeKNG8OPRh8pA8+vR4KFFU3qBRTKf6K4eQFqqqkotgTYmomO7+y9ma+o3VMohxIPJ4/AzjtUa
ebXetYTDODsp22oABtx1jO7tgQqInlTF9TidM8PQXaz587aWcD2uE6qoGlwFRCj6UwBNbiy/kFR+
IgpXgoMSgt39n9fBEhWcrAK6J/b/4TNwp6dEW75Bh3Gm4Bt8lNw35MxU/GQ3IGK6UmJVbwuixyva
wj4SRAzL9MQBcfbmErj4HuUFq6+1QEMmqMZyfEauuV1EFt8JNSxGYRtirfcj+8v/SuRe/JVQUSd9
Dug6PdCXfoqjNapT/5C0MeeOc4ycxJikiNoAhrk/iQEtrlV4oumy4mvRbphopwsCwU9LjWP06GlP
+t/t/3692QsR1hPmTDVI2gjtlbsVmfkB7cglmc9ss56dfPq5jh8brviUQSkFvYFWKUF7Fk4zB94h
ksac2ywqKCSRgzQLhBuTKPc1ykTeZeU1bouKDZ5MWg2TsthCO2UYcI5HLKJ9WX01ErT0Xj5js9pB
0x4KWmkaPPyvyGZuDzZu3v7nbZsp/Yt9h6UrVnDIR9BBW/hWFSceXZMbHjFPLkxuRmoNAjHWj4cl
S4ZgIuZiFjE8Lmrlw9slFydH+CfRCZZksMFpFIPe2G6bNpj0sw4FTflwBiHbCMnKPp4WB5o0DuFv
HYeI/dQcdVEdTwJiesLmTM1Xf7GqAnMGl8bjWQ8vRyvVlb+b8ochkCWmRZwROPM8aWfNJEp9iWK8
gMYUUJ8OGR9ael8yGQKVzmH24Yp/8HzcywnwKhfM4MRJrYoX6/Sd1xhNysGKBpVOX087ljjspqyE
/Dpe+ikTStQACHuq7wZ4se4WPGkyqnAHZlfvOfHAe0Kh3pqwdXJ0enl0ML80YqlYBobAGkDNFYu5
NRU5Bt9QUuOSqXOMwlsTy0wdRmPyfZdpx08lYStTigsoFrCm5R5de5gIsgWTeL7/fuolZYyDuxTH
YswCKW+mcgWyOEnDZcHFI1JT22owy2GyZ/+06NxIM2gm0RCKOWG7C8BVYGCR9j9d5QM+J3/Ze3f6
5NO5KNij2TQ+nNbr/jH2hp91XIa5pY4j0w3j9MfretC5LcRoYAARQIdzMind4xk0zATElux5rNbX
S0rCdoCVrTSIaSRNTxIjQSPUOgFbr/NKGkvOupDg8Kgcc9x7zLmf9u+Zk3D6ZXYJB0nQDqBT4Wea
YDOCrrzmbfPvlREMMsOGJu8t61RzX7F4vbHDMQsqy6g9qfoybRcAhiBYl5z8AUGeDxXkOd8ztdnV
fGjjFmJGkzgJbiFPwMWzJC/rwXr5iUmhuT728S3JyN5lQsmrZAlVV13hk13VdJ6+S0jUliVHatyc
K3JwO4C7TABbglJGYyaacPx1Lg5UXU969NbFPo63jM1eZgqywDoUPGmgAhcP2TN5NYecCpEiYzKb
6xvxylvXInwIK72dVCTUaHrM0pms8+ONPJHfOuSaJk0ZjZeS9rl5+5wFuH80bN2zhkJtvKP9bddr
HDxHtHloT3sr0pWNCWbJ0FrdRoFPezrNMduRAoAjfEFUf0xpi1Bm/f6PwT6Tbl1ILTI2erPWRmoY
gfqbYvdN73mIczsrzC6JkdQSBdwMDdnf+XZeSZk7La+qMVx1MtWAwAjRAehkPCi2+MiyXTqga2VK
IoV2pARuvpdbNPguRHjdx9VS0gIdQuilVOXOGNWtedRQaS7xjuMvodgFYQ+41F7/UwL4ONhaa4bH
aV5xdmD9YLRthyaRNqPGklLO6nY4QhRT472MYxq9sm3L35I3rgkIUI2GXW8wwKo01fB5jEqd7wu2
bup5MDkcmmfu6SpbQq7GGYHpjodLb5STaDOj1cEDOCv0Rp5NpastT0daVIEDJU20JKxlYC5uKrWV
AABPd0pQ2WzxukzwLIvZfAUj1uHuflFRUsfdKVV4PV2JX5D058jfNwpMYdhk+04a77NhhoWOfLX0
7E+vaWJrSmHQKnUyiN1V1MGGt0+iqh/8+s36/oG/ZaaKM07Y6UALm3b7wSKguDseatTGQxIlALWx
GhtN9w+ZdQevnG4YDR80/hlqDIGw9nNX1vm4OxPmviBHx2ZeSr4OnH2hKVEzy70vIk6ivS1sF4Ls
/iaTfwNUEx9sBxVPHKR4Pg+bKRhrY94BfRMiWSCHzRM/T6J9vY0mqXNEn5Bwpv8HAH82ZSGWCcNt
t3lB3qPYFwB9WNujUgAY8d7lHBD6Jnd2psH7CNFKzoYdZDyogzTPdJmOg6NGAWtlK6igtd/AyMzY
UuBGjWEC8ScxSLDhtbOlqrNg4fNNVWGzlV/dCGmm7GmQneslOLAOGtH8vmMBXpJjjM0mqU/8UkNu
bjdEuYYK14Pjqiwx2zu05wmj9qTb7HYhsE6JllZTDO0/mUMpWjhwqYSCgF/bIFl+N9uG4cOE6Igt
4x56gJVpbFMCr9H54CVdZolKM2QJ4dAfX6dV0NnY2+pudFi4cVf+1CGxa2tf4Gc0WI1X/HLHiU3X
xfncTLFbKFJuQWi008HWoHdZ7aSQ3/v9dH59DRmPiF3Osu6pLtXyc+SVOLV5AfIRwEoYEhouZpie
69q8vPbpve8yMzasUBQgWTZA0kF+6QXI8XlrhprPH5slKbiTsy55Fd8IRuVuBszFJoFYH4cbRor5
3CzAcwK1BLUSsk+NxyGCZYe8p3ePgQAK7W1DvNKlqIox4ixqh6ZPY5DZ084vNwGqEyyGV8kXtzYL
loSTxNPRduc0uBbN0nsvVos2jmn5R0ScubkE3/V97kvAr/JQ/iErKTCX02poz3UKt4TjsdoUWXyH
W71o6/hTZ3HqGhTzHLG6bBMC1RIgAlJgFs8uloX9YiNV2rOWoN8OK8pe97mqaZFUOWhe+mqVLEj6
QFXjyHeHRmY0pewkXgN+7gJN6X2UDu0nXEmo2aS0FKYW6F+ihc7YEU512GlBxBHi1gOUHYRGrc6l
0mtsP1Wm0Srg7FRH3oXyIMEmoe0EgA6gj1sDz65J/BF1/u4QlPtRTpkx3aHnd1IBDq/tJHFUmnWs
/kyIBTPt5AtB8qr7QIdicxSaQDmHXPjjG9I4ao6kFkJj/LSS5wEtAHjxuh2y8M/fj1zOx71Xhe00
02g8NYNs81svf8yDsxue/SusZ7P08wJ2xMXtZX/cn8nz0Nemv1voUl5yiZ3a3JhTapzMGcNTfrgY
OpdcXSVglhAmxAgwpu8iHG5OSaeosztVUhTMAtz24A3g6ndf1gz6j8sHuuFGLewU+ySbFwUUxpIV
q8DFpZPzxbOh/fQmF7M8O+mqgIV+3VqYqXU4hd+B89mq36FHUmdnTzOucFUCNJplGVXbUqyaq4Rw
C3Fvj4Pocg8We0t+xdykUcfj4JSf5mCFF1FvCA3mK0cB4Cf/QRTTXR3odg9pbGLQnWmUvbgq2PFw
eQjOVz4/PZT1iiTJjsxvEr88PcDnlVOzPEirctOWT9AdIRIplzU/T9SdD4ND12OeHQUsKlAMoDTh
LHw/3Nhs3T3iTQ7JVwMXynfGUL5cf3sQrzdBoxBS4t8+9gF8KcJ5UK8dtEKsSX1VR/2nawuSjFO8
uiOFuhvyrtrmClkj+uigcLs6DmX6C6WB97dx8yc7WbDWTymA53f1h2aorkT3oRhMLZdxV0qHALcW
ya7rkMEe7QHQ0vscdELDW7SyYtiXV95veN5m2lfrCoNC4HV8dvYnmOIWonrpIQSPGYHqNoJ7aD37
zEHK/lNW8MKZGj5uOMUo1OsRP5Ynxu9CrdrMMO9sbEDJ2Yiq58/G2VwcaPwm/re9wnXXg2lBGUsx
4YVsvTPbzM2av0g9M4ThqMCXoJnKAcZ6PmVbnJU/ylr8B3r16c3iAqP4xOdM7YaUDTv2uFG9972Q
C0qJ8UZ0BlpjR26rRHT2jlyzFBeVaI7TuDaq3UxDmhaRjYg5l7A3I3y+Xt6xx2XYKJ3ifCHZ+dA4
/+ZyPVRvcpnwsB4FVhfjJkLHQLIpOhRwm/4mBGrxJDJVbHCPxxx76LSL2zbWZ9NoVLbV1MNO30zL
SrtU8pe4IuAC8MUClrMEacAePcob5xn6OjD+iYlaPuv5SEdK8SSyBVTvzBFOhXx+4APWp5Zmeiek
xMWxF5S75asgxdn44udm8iJLlTW8CIAdRqbntc+4LSUaJ7DsjnZWzzk8xq332Tig/IuA/LdVNCL5
pyVwmN0PxPwUgwGEPwotFdXlyirSW2Rl2w/Q73qAFvPCl6o8BtpKtc1TIxM+kz7oWBT1eME9sRS6
seaer7ONCOEXHDR7zPCs+c2uacQkJEv+5OhMudsckAWqdkqxkevlHC4UbGiwxFDwu1GmnCwAcYxt
DkrHXi4z3qt3HS0NlKT19R66bCWH7jGTp3kX4fr0e9WK5pzWUoXbMyux79QP/BGsuYR8tkQeUAPY
s42ArYmbuoF8SiC/m1CLE6XVqEYPKpXOm3x7rzpYLLqDPxE/seR++cR/qOn/Ltfjmte4YPSCm3jH
F6v+5l8pVYnb0p+zQHU31nlm47k5jLVXmbznK2e+I3FYjQDO1jVgv3wvtFGBx1ZbibzI3NJrqa4O
Wm1zIG5xcvx3uNtv3CIACwGxD3FMS57XnE7EumArHzYIFz0HW7XGC6EayUj5L3tlEa3Zg9aTO1eU
LdXalsikhlb9L9LzKc95w2EyL1NOgwMNFUvMZV98glQPxMz7UennNZ/mt1KhOWhXfAKPaHEwPL8M
+GI8Bq149NufSsC22gvd/wC3x5agtNwpc+ca2vEJT0qLjGKmGGMYwX2tRXXIXwZMBMITQKRsnzs8
8UDhTHzhL5BWuMU+sIljT2+Pfx+Q7RhHt7PS0HFXuN7kG0klae5wrJhS0D0YfbdlX/tfzkRPSF4h
P6ZV4Y/CR6rg8D9IC7QM6xqJcW089nfFCYnj/WclrU8He565ic13+yv0hx1VdQi8A24Xcs69qLFi
4GHX3Y3p3EeXTbYifGm4ZE6RdLxN5nvvCcFUUT9FexJksxcL0qzEBfMdakramo3OCAZZ4juEbQdo
3whf8WwJmEUr7UUTDczyOIONwcrrdKWiz9EPJ+CCGbR8BTlZOY368zC3daZEbOkgZTJPH01ivVyS
ZLL6A1yNynYTZUN8wG/Z69RWJdi6smQCFJNxYwUdXCFNPfZRtaj9ET0uLrTjp0/onl/3JG5DizxP
uEbIjt1giDi6wGlPe8D+79AoYTL0a5TaxxbB66cr99MaY2B569oGIsD6qUr/p3cZCg+gtk7lDzlt
46T7l11bz7m3u1pwlHZtEySri/y7gTVciM9gZZ/rGQi6Pu9L2tGiJYrjLuyaHfs4y+VIycWPIx0F
BErq/YnuyanaDEeI18r1ONIcZSqy8ZFdxH/uuub9zjQQ/d/kiG8l4Xz30HYCS8Pf1q4I798rcNxI
4xVgeSOIVJKiLyjNd2oaoazV5Fda6PrvArGcEA33dcU+wwQ5zOJBRP7Id8/BMBzT9R0Ki+n0QP5v
IR0eJOtB7WucpDJQcMQOAJzlGa8XfSmT1Q5GqhyA4zt59euthh767HoMKBnwFBudWuUzC6wd6KWO
cqeIvYemGAJ9j021OnlDr2F1P51HfWaNeFciRyeq3NntnOF+Q2vCiaWjyDIp84M8fhEaqheTSrYP
mnmIqDx1oszdMoLKPL1dcbvBhrNxbspMJPPSugrtyYN1IIwirrFXdkgCHmDrEDbuctLFIcUA4CcY
FvpDhygyKyiuER+ou81xOocJY7wUcFX4Vvkn75vMKfLj1aZi8BxoU+PK9rIs48kF2cUOpyvrEgGC
wbpgCDPmZ64zOtWvuRY+B7sPfBVoIkmfDR/Vp9v9Br59WZuMQep69lHudhci86v1LIIton3aUsLZ
NZwX7CYJ+syczqbpgMp0OEK7q5Tdc5fe8lHm6rQzwQUAE463t6QBmc6IZkNSRbwK9IwiKq2oMZc0
TSeuHOVxE0x+AO5YGtEHmkhbJCSW6v/mQVAeUSNsXeH+5p/uCc4TfmkaZ7wB6EfUrCgc5gqWuDXx
1U/gPnvk3jF4mn9vi+ElkDmi7ggsYrVnRjXVaszzC9XveOZW8UiU2cThSy752QzmCDghQpXdVzcP
+F3hYtQ4IUKm+T1SuZD8VJi4sA0cPJw1Dfmj7HuU7OZvnoD0TJytnMbOdQnRPuqEMkQVGI1s8uUK
RW5lqFyaxHFgMg/Eq2c3p5RZYpvTnkMNQfIsFzWCPYpF78kOtQjBwHwOxoW12zXuj5LVSJ+meG/z
iJW2xaadWnAikKU7g5FbuxWQOT17Fnj76mQZT2ZNCPVIxtQCVioiqWWfFVPW/7hL4RwGRVqpo6RP
MaaT5r13swVIi0KYhd3mWuXf9C1LVBpfRNolGn8O+9bfKRQzXLeVC1AnOEAUNgiaxeWXJmQtRmPd
XLVRgFUbAYjJ7HNteV+fZxwYW7hdNhYwil0lAlj1yUNc+PIBUIkDzTEx++9ceroQBJEFfNp76OmN
Q8oRg0sTcmnIKKgXYm2cFIcLXp9Q5b3CRiCN6fFhv0Ko6EDOt97xr5PgRlac7zq7ZbHERjs90BsA
3ZbVVGh4Ljw1HrAeQGd4xSRHWP1vRPNPRM+M0jMt4Rj2NsCu9nd0DTJDpqVMi+eZSiWJpR0wLahh
0q1z2tpwq8jyZhofQtLAPJGbs5sTBwK0bTeEbzqqj7NWN7MQ6UNl1G3uWdRP5CLBQOniWcCBb7za
RCO2Bjx934LPrVyGEq+o1jJGiZUSOIUp8mpVQEYw74Xl8sCgLbtBOjdTcjIWEZO3zp1EGV6Tqcax
tJ0uQt1cyyIDlP4lR26NDQKQaSlle4z8DJ4x0jzk87gQckPLLU6LKNYNSmt/0oF9abrs3gaXa/HX
NOvJ4NNih5ViPtFz8VlGG2DWvy6TKERvTOWD6JnMLFC0bpwBBypkU37Mt4HYXxSnXvRIPHQorys1
+4piCn0TgHX44yERTTB4IrBaG5Obta8U5PgdlsmlhlXWkRPL9wOtJGE4SDx38Z07p++UDYrIcc+4
5JWNnSYzdBfsIhw2f8gDN+ljF4rAA5qbhZOqDVfDIZDQH/bIDI9SQHa76zxEB63dTqzffLYx17kR
c4J8denVIiA7z37aA+AUsnnKQ+Vw0Hi9M3z0cQTFp2Kz+V6f2JMdUBnYcw5vkkzx1oaUi2ptn8G3
NyJ7To7OI2ew++0WyJTCW3hLtNq1gn/gS2/AFkrRrtGC1J9oabHo4sbOoaADkEY+pgytiTE+F2Uq
moFZOhYnBQ/5lVmkx8B+2rQvr7t4vJcjzRoy9bx7MI3i7PcHioje/FQltM6bvlhPGIpGIo1DSN1r
hCun7WLxnHSTVvY7bdL505/ciY6dO3K6xR9F1BG3RhYg7bFPgC0aezS3tWZptMEkWUziLTQwHIcq
WJTDALnyoW8y0mRbBnXYBV558W8rhy22O4Qr9Eawtt7x4IySAqln53aHxQFFjCjZfaMrvv5BemfM
HJpFoMpFm6KIywmqFT7Kt2dqDBkcWD7G++wPGoMhkw7d2uI5/HOnSZnAjbxJHcqnRgo46cz7kjyz
EVT/nUeUAnN/4VXAWtTGwciauHCstm3r4oUrdhJu3TyO4ijt2fbrwQ6Xfrlos7JDgve7IaxC5AJT
ic4vTRiw9uJsXnmtuXiOwwl4rxqIw5h/smAW03PxSfePnXEdr45kIfr43hC9Ap2PZ+sHYRJL77/w
FMyn+hkSFUh6zhtTVM8QTgqJBT3gZiaKaZn6sy1KOyaDeF8lH4z3g1kHbGxhtDGmCOWH+injmUIN
IrH/iuY5KLk9q01ixKPqGy+CsAUlKJJr+aEIPyflwYYzXZPjtCuGMVAeS6ryTvJ2FswAZ+uT8ypV
KY3Sqq65gazr6Febn0oBEsxPVRknrUtFTVCpChNqKgZ/rYYvgC9N/hkjS5v8QX+zQ9b/QbHn2mNF
7v/GE0hbpFaKXK8QC8gATKC7xw372T6hji05JUPhz1CtBInrkR+v/FJdfAjtL0EIxRQU19gSgzD9
q/L4ScAtrRGB2Q14T/r1LlTlAIWqQNiu3+613UFZSvpzwa4+3r0M+2ndbuQvV9lRxaKL9nzUXayj
WqJWWgqJTt6veXORPwjuceOI3VROE899ia3sVeiYxyY45uXelZenw2P3iyc6dIGr1vTy698ZOwLq
+Tj52H7ai9IUyo+Ouz2CaaOQNWEqJSVbSWD8cGJ+ru38CtHQy/yBcwD5wD+Z9FaUGAxh/plC40sF
8n2/4kENw+ZERcLNkPFsO3GYKIthm8lKHBC6MBJGHBg40lNebNnHhVB5JOUwr4ckdbr6TOwdkq9P
EKzqhWdChveQo9p3aD8rQfPmUkngfbE41JuHBmAzZM8eAInIU1ZytfMkMe+qZh9BpUEvCcBUdIMR
NIwMxR44xOWxeXmXc1TRvvuYyCDefUiqQLgHip59KrjzgozHZKHiG+RHWj+yj9WdUbIKmGV0jwAk
m0tdKUTcktjpIahxM3fu08Jk9Oq6fgWDDrPNYdyWEUDHFv04PsE7vap69yCi4OaX1bKog9yk3DwN
W0idIU5Y+SXz9jDe231aQuDmDWs8+y8hXseBmr1oiTfqJ6FaxLoYS9JXSsO1sM3D7pWrpppac9fJ
2zFc2uOA41fJnVZ/4kUfM1Pm1G82uRkx0DhA0CIWWg1W9DFfwixQwcckiAEAZNozSE3EGJb3FOlA
9nWjWwd6+gE/7T7B+aaFx+Le48PnXEPZNSNao34S2USszTMRIkU2kZouO716/AGeZSww76mAYghi
KERKuwS0neIkCXCQNHIWQjXWGovUGiEVwWcfTvneFHyx/gkBQz1b/OC3DjqvrwGhId1ypgawjyte
lQ3D3QN88vzQhYV58PR7vKidDoGQBoy0cn9mrudmHZ2PPZELe4nl++mXXToSk2WCpWR1c2Zo784/
Y0l/m3ydFIXD3JZ17PxZmgv6o4zOqd8kLR4YJMof2krSG+TAjbhtK7/fgozDWYQbjCvOUAHNb5yA
LC8noY/RJ+GXLRHUMMfQRSc3fVTMre3N9+S1ajf0Qh5yvswJVJuqvfddWyMdyco6DWWjyG0AJZ8J
f/odp0rjiW3yU2J9pu0sLfHqWFbK5aliBl4pBMXiVU+ljYDRQBwf9sa9DluDDvmj15kIEwK+gn5Y
GzXJWLLru44zKh7qBMyYdltXNQzxswt5tSNArmaROO40hfVrgMbK4xZFvDzNcXe0C7F09iaoybkN
jeIeLCkH4PULV/BFcJAA9gEAns9WQCmu829IlhgESJ8HVrlBkgD/f9aqsci/jsN2xkqX/QDzdtiZ
cMO8swjrDJ11C1W5b4bTeG17NNAEHaGXdJJ1h+LG3ouenUibjfMSuedN0qZngSTVca2CMQVKiYD/
kJ8te2VLpzSc4lvUGaNViphlIHSwvZ9pko1/7uR9aB+2/fOKdGJhp0/1+Rzy6UrhAfVDQ3I/A83O
TUtohKy6EAkGL1U3ImKmOcZ2fIyMtJZTgMba7uW0vRVqXsJMKEaZTyvW1PApZ38aZf1RsBb4/nNZ
gAdKjszbfSPe+6Su4ZcO1uCd8F2NB6NzTGVvlpz4WiuXi2n70rMlDpQMKz++X6SRKwESURSoUPgz
xerbvlK1V3OWK2YEW6Qo6i2Pc9bIx9mTnUP5kuZwVevt4MnKjc482eZTgvmY4VnPVVjtgKnTJCHI
3kfX8n2ip3B5gIavoGHyL5elhCq23GwRqH+Yb+yEbhlSko4s73q7jTIS4cJ1DnUM5qDjF2vxvTjx
6gIgmuaaNYV3xFLB4e4AVTve7Pi1j1VjoObyTJugxQnZLHXepe6AVwDKbHxSHMyy9D2DUFP82RKs
wHx+CkD7mwAir/YP301FBGR7dG3ou7zZvgKgPm3AJozNlYEJgafTbDgpufmN3y+NxdDRgAK09tJt
ZFxk5l9AV8ThiKJhQYRDMzlBo3KdTFvPjHlwUWX1vrqvS+CWzx0mv9gMUN/EynDn/Hg622v3AWH0
YfS8bdOyyfaJfoJAGyGP5sp1Usp31I+TMGcEkUqsCYnGV1yD5//f1AgelZfrBGLUrvdrr+pmWJPD
6A2WIh5lCj0PiVnpNhkmSW/gfj42QCKmhyEeg373b/fHkarMTQ7voe80asUBrXsYB80lyccO38Bf
mGHl+9y0dxVD1x2SYM0tn+j8Rzn6I6SDmXmef7ALBB6dz+oD0SO4Ny+GJoRb6jIMRXtIEi245iyp
61wpcO8+r6KLKW/wsegwNftYY2gkYbF4ZS+tvhhMOOSf5fLW55KmJmdnrkTDiy/So402wQhVwEi/
8Q7aYFhJcVYUXVPik72d1/QJobghmhJbweZpKYrpmiU0W0kMKsscHUtSxJklTsvkDbVV2sA9oBL6
6UFh+1d+UghICkv2YxjzUcNKOnHj4PVwhHzCEgjhdAL5MOy76jiZJHHWzsFOHX6ZFdlNIsE+4Xcs
OQSSuhPTbp5y1GhLCv/eA8uBJvfQ5MqF+dSUP/AOOEEYVL6TLRiqGpx2GHvvhvrX/2S+KO327xjz
bZ5htc3Vg0zJ3pcSRcywtSzwFTQdZUeizoucVsz8lMRFudS220QFKDoP3dfTRvgC7MGjKDgtUST3
6l9UsgCferfxXX2Gb24LZsLdTS9ijRVnhkQ15sbzLE7lwNv0kIxTzd16m6HZfaclTz3jxtAlLs4Z
4FbmxOWf9AuEqzjoL5+adyq8KJN+YSog3MEYqB9xReW5PLBeo1mwKP+IpFLOwmwPOVtxYSVN0cD0
lCOLDEnbBMLGHNselXtPQKB5OBDOJptpjXwAANn/brsfIZYyPWs5APhTYim0rX0P+u6xiYqy+POF
+Ec9MwaA2Enr7zxAemaN+Qy4Iqhti/Pe37OubAsKu0Bvue9Kxup7zvBONBbEnOv4XM+bID2uSKA4
kYgdmF0LGMV1gTnG2G8ZsM55nM8e43oqCtDLEaIwsoyifazapxzYMmfJYDAu65jdvdjuDl+XIj+d
izK5eXp2I1MtxO/3nMrtLF79455k2URr2cGm5EDwCZmCAVO+N5ky7nN2cTb12snV/Cdo7enmbn7v
0t6QGapf60eZcS25bfzraJO/9mlsvTTk8xBnmq73LR0Gt9XtE8WU7whcExtdbVjxTfr5j8ke6BL8
0i1Hq/BodAwrL2zjT4Sj0DJOSQKKbGRfbbE27MUMLvdifwKiYz47n5uE0MM2GSQMOR4NUKbvV0PE
VMH9ySg+ncbXn8jUGWzwjcHwisFYJQzmG7/UnJHja0rm8F3RgX+xr16Se8JM+rekFAajqqa/eAp9
/+7mVTHc9WTeCggN28nANHypNYRIGf4xbBQpiUa+iC5TTEmbwvFe4XOZiE/1uKX74+Q6CgPOhAd4
2ULdnuo7v+VfTri8ramlrsPRE1KVX3EpcG2GoJzfHRCbbef9d8HUxwRKMWSc1n/rjvsjr27EBd7V
F75uMvCIHDsxVmgjGqfInCFQH1efLVoM9wqtFkSlP76YZZA8lYSfk+MEx2PE4RxiWcedeGGVgi2I
P9fME0guJ5JQbjQw6U+6hUWLoq7cf9fNXac1zl4A76o7pyMRKaIcl4UIhbdp6iTekmvc1uJBd9bs
CwX4RUQb7x9xkOeWOf24T3Nf1PeQCoYEu/tW805Wj2HAahb/LtPlT5Rwreo6Y6Q53FWf1oUy/RWY
GeM0KqsGX02ch9OboeEkZ/refMB4OeCSfTfnKnlEZsmJTkib+hivEAxVDFfu0EFzSjNUdfm+R51s
0tdmFp25PEg5mcrop1fARDns0Ynh88/rhuRWlLaTwhuaotK49Z+58FLn4W2PoHkWJr1IOV+v38Dq
M/CWP+c5+TAUZypva8YH2++7Z/LieI+aI68U/x3kJQYyNnzLWzcLpbovGKaPiqecYZF4mQ0c8n/x
b6oSeN3Rai+r83GMXu5enc2th2c+sMKmcOLtK9c2jRr+swBPe2y3MppvTUSlgA9p5MxJ16coQ8y0
A65jhOsEdqmcSYoEVxAWdhm9VmrHFHbzHNA8tCBmb+fO2NWXY7Fz4HGyw/a9GLN4pNIJ7iRqcSTm
EG5R1pYJ8eI5MoxKbwG+VIqYTksvfYZWP/963E8QLMmzYC82w9yWXdwGcv4WAJdIe93+vV+Q61Tl
eIGHHg32PqIcXgZWFrVvTFLZGlXE8Fc6j/YbiSz8J00uQ//QCWpKIY6DMSvcreOI4USTTRA0uHpy
6X37Z+eozNaPGFXp/HXooZF4PMLhYuW6KuYvq31S7Ojuk7V891AgJvfncjL99d4D6PwYXBMhAAxS
spXUEapANpNGTBAfP9ZDqP3IdDBNSwc21Q70ua3pkZcnCD2a5uJh0sf4I+tyNu0Lpf68HyrqxiTP
d+ylnMRrp97WmR8WhL6EummDf8dmYbBfAOSzt+/oK/lJkq4MvR1U89Mh9r9Fa486i/drVsHBPD0t
nlCi07pSTtF2Ei/+MF/nugri7sTveY/A4Cq+XdpK13FTAVCU76TC48/QIU6e01648ARXLR1jR4rH
cwsLx9syF6Tid1dvyU8t8BuHIGYoBz5DlITV0sy4UlDCSQ/UESuXq0DWYi6Xms58igpARQkYvtFJ
WeXC2qNb4VW8T3R1SQxVPB/19uXwJrFhtBLaCUS3P7venz2ID3pVGtz2zbrYFU7SOj61h510TxTE
fkOcyIaOmQalgFORLQQMwGw6kH+Pz+i+PZJaIcLFpleRJIAXK/usQvo6B5WliB2of4RhvIs6ufNW
B/PIqH5m1yHgS7sgWsF1JLIduNdigV54FIj/eWcTQW0RAxh99XSrJZtVpIplld8UbmU5pk8ogx12
tQ6wOg5ce7E7Y8+lNhwNAbz6tSiD0+O2GtvAW3GMlSI3mnTBTAsFTTY4hoJehfn9oybK9twqwTuc
IUN0bGCRnfpSvcOQTPdOtyHlBB7E4bDLpMtcCHlI3LU/b9Ah2oD/NFGsf3m1g4xQmgXr2MVGIQ5F
a5xB0dF51LTUNkSIc1IAOGzUEc2vdEyMVswPwKV1W2laGuwue5cAi2OPv/+mPswLx/bH1E12lnzf
yEhBi0IyDNR/d0vaVW7RoUinsTP61tMPY0VVGpxg8d/pqC2MV21lt55ckWanwXttWhZxPVqwry7W
Un/z7YjpOc1ANQ0GCCWob7R51PS0QYauM8TRc0WNL1emyYm2M2pyrOeyy6+EwcSmCNPglF7gWGCR
dDAJFWT0rsTm1lyJYo6fPtdUhm9eDmlRFST9QeX/SKokfykhTs//k3nPuafTon0W8Az5GYI3zHmx
L/VL8S7eDw5Qrw2XEIcxZG6OIJZs8kulmjYlh8nE3+LkMBOq2q4Mj/4wiYSpwiGaFan0uwPdLRpO
S1IBh869P+ljE3XSCvf6r2aprpR6rpA3X6F22RksBlZ91ZDHq6suo+dxGIuoaAd19qilANXgYQ+u
6WJzUXblQme0pml8dVwg/3xYMj+SB2C892j3jabaZX1z+q15qLdXxGBjrfRBbMrtQ+76Hc8zZbHQ
MfyUh4cJI1gcErHfXRyWYxKI2xLaSeVCNPWhmlElEm1wobSMhtYuTKHSxh9+jJWVIJcFZaP5vx0w
HSiocLCJklz0MScVU5Mdet/22La41oJPiVG+GY2rjFQYTKN+oJyof4pxzqH7vkUllMNwU0mPRIN8
Ctvkl/sCY84hYm2xviTCVBhVK03fitoEYIN8AvuJddaGErz8xJSUFm95uWu8/9z3LW0SlXy2GJUo
zXw4MbDdsLtAtmZ5MK7RxBRm535OVlDAyetxFuR5hPOSFISx+X4YqMy/6yEjZzH6nCVgHvic71ZJ
Q6eqLYvRQpYwmFckJDpB2kKS+xYjASlxReBQAXuY1NgPe02lDRt2iGOdgclOcWNQcjciI+kF9GJA
9kGHza4XWotgK6xpusyGccM8/npsMB3Q0tCOHrs7SS6j7peGeQb5A2lpKSt5JYTdQbEj9g7gneJr
0FYEMba6RPpTlEXU7pZJbBcCBwMpTPg1hwXjw7M8P13wpQ+cK/vCseBw7AMlmHasdjl8YP+nacff
hbQFyfgdami0uQIh1ZROrvKoBh7P4ZIS3Clk4IPsu4nZqeIOVBGH5rGsk/V58vagWdVPeYwed3Rp
S5iBStF1oEW6YZUX0q+MHSgc8Tc513Fls31eowTJDUTXk/Zq+CA28vyZ6Lq3N/spdDtWHrd6aATN
Qoi+j4IFn7mMyAR+UipXMUqBPTGT9TnyTq9pnlyO7pSxLEGK7u6c2UYpxaJzXeFLui9iqQrJ3VSd
RpsonhHisYbwk9PrMaQGm8ZoADG2TWPOHVdRukgjALb3a1XUOWAjN2glgV2Sz79OhEdJaF9VjjdN
nVjam98PCljy8Pr7z6Ba9DjY7D3FIjSHGsKkPA/BEQE320Ss1JmDhun0IyY0rmYJRL1jf+7Jz4Lg
lYM8ODgD5uVU2Sn86Mh0/yj5P6HJruCeFbZIR3z0ORQTJTikRHO4jAVZHJ1qTbNPXKEd04tqoHUS
1BgCur/xC442ptB6VULaBt+rjQzHZTYp6g1+8V3cv0cIXcx1F/vVEVyGApyZYav0jImU/A6VfnaT
kkZED0FOX7iXSk5ZnirWfpkgAODPCkrS617U49I04ptfMqXV+yKUpB41CVDYYPKp8WktddPo+fx+
dCK2fP2SpbfaWW0hyGkCyZ0s6asNIvUgDXrUYX9Qq7jpHvJo1lN+HGvofigZ5NMG0HG8nxUTP7bR
clmm2mbfPpWLfA3xtJMvlD96bsWrxGh9cJq6r5B/tbe0twFAz9c6ZI6mS9uZEtnbRdbXRkXimemv
pst8AsXG8/MVIZuXieBdkpkRh+iEBG7LGnJo8w4IXgMUZKaF0by1Qxtg1SATLAECxojLWmNtyB4G
f5npVuboNCqwsQ4lSP36PYrpD2uior347X9wdafJKfByLMUJhUjbxWhTnd/mJ++a1dz8QWIGoi6c
Wzld0qyRLadiSl19+TlVbPBSTvp6H+3XfLMEFL1Smy3dNAykB7dIUKeAACYy5ZogfumcPnNV/wkH
xfb3vv/nirBavAz14erEKRyIlWaRVC5dgwkP8FESE/SPcezdQmoCVRhosDFIa4jgCMfX+CVaq1ir
qCb6ZEKRos/5Xu+w4bnntnPUkZdfYyhFUVCBM4WL/R283wfmkHDb7UWpp5Iej08iCGEc95gQvAii
S+gsq9ohy6wSzJUrpFbse3NPHJURHl581tzLEntuMp99wnCO7sSGsbN3AkvmRPGgrfbNdEEgMt5+
cARoaJG1xDHdV2ZDkwD2WLcv95rOKMNCKuR22TtL6A6BoY77V11BjqyGyfHVd9Alhki/nZWqMqmd
9h5A/ujL+8HTnCvds/C2sKUBkiEUosZDnDS7sNNhdDqMdyhGv1jZYP9BeaIMJVdS8Zw+jP9hGMgf
2q5fHoBQ30Z1hZCmQlQjlvT8ce1i3WHMMZOSn1zm6LMawwIVmceSbJi1u/u8dWLg8Shw3B6wpgQo
P4u82jxDJZupC7s1rjepzeQRFHO+lA1yjWjZmVcdpdogpbbCNmpRdnGv+32gYuHklLhhNr5iF+nr
otgsY13FR0dwe4PGDxNjgjnPWnxdy4pNFOeOVV9qqLtElcY879dxclLP6et1/77hVVaD+dhwVDQN
gH4RwCYLEC9zf0ZoG+AmfXqORWqVdgZ4P8718uAbu1cUpjWE4BgMuOy0Q0G93TwkkOgq3JpJBJNS
xmUuGXft+e0osG8AcaQ583JKWtJe7aDCO0FXne4D9PIvRAUPIrOlSWEjZ+P3RMktnyoNIghN4PYL
xgFA5IgpctjJwllRe6lVgvdtKdtl4FETsVQK68UZTfIMEJuryZ2q2OsFF/pPEq7b5Vwqzb9r/V3f
b6gOs9V14oGUMw8RemT1kIIxvinrXxMkeQXo2NYWRIIoYaurzyqnZJDbY2TAf2WJoG5aEWqZ9J7G
0GbxGGk3rXP9H9dDMlvK56cCNRCGgGl2HgZkdcN1qTxYZ0Ky3a0poxZCfsNK7sNaJ3nOw8wzPH4e
ymtX7sAmPJ1GWVjIoRkp9yfGIaMqo1axMdVMjQICMtlOyT9+8ICf4HR8ktg/AV113uCxHnZw7SKz
GMEUk2VCVHZSJaJ+SWofqUFxa89ZtXHnxoPup7IqCpQe9I4sZFxR5FOzrkI+cWlehX5q4d7we9CL
jacXQbJ+udtSNwbWtCTLimp8Qx3MObwnBbkmaI4JYN+tbUbvZqMxY6JVViHb2wDesO6GpjDRTK1N
P2BWJirt40gNRCAFDJsCxpcXQeImLDyNankm1AVH4nOdX8VyMDT4MY4e7tSeNCG5e7JLawTzNl22
TZ4mu1jAgkm6y47j5C+UYUrrtCspdCLTOmZy/Y8glMNZvKwT3vHsEY/7C44GrmplQqgdmUVoq86i
40NfEdfN6+J6ngBTHmFV5xj8iKW627vgICEo99hpm5ASjHcsVzXVKfUk50TWwy7kQfo6X10oFHjC
VDjlfTFdK/KEDDaIOTWynMecZWWMBKiT+WPwpT1ZwUMG6l24WkdHNrcOmooDJVI/9cC62oMHVwXr
tBtiWG+AGGoti4KvNlMJS0R3ScaF09mqvkbwZ6DgZhVewTmYqZ/bgsU7/Es6uPz8kjQnescQi1e5
vDSNEnImVPGz/6ynS4TeQdDJfYavvQEN32OZM6B52wxIj+/oyAa5hgd3Rr/YlTOXg0aplj8fFsE0
grAswnJXTWMT0UZ1yxVYdutGJAugURdAo+WKMHOwT75Xmk53DiuFRvDw129Jta5g8Hs+gJzuw+/U
+uvZaysSxHmvXoZvjY+b6atPdPzikgVtloQdu4K90pr5MR6/fZ+KvTU3XmJeC01H0510v39Zj0An
Dc/bIU3gbz3Wwg34mz6czXfU3qDL1S/1SwJu4TGFMThNIITxvZqYV+uL3oAxB07mKFSsq29FmOb1
MYqWfBVoNo3Yeyy50DN+Ws8DQHdAnQybHyFbsQqR8OHNfRjknUBfhKdeCBVglzyrO4NJRrnzb1tP
h7ojg7jTqlN5Sa9EJPoiHdgMg/JA6vdbIH4DZurwuhDST8PMStynSZuhZOrnWOsInGS9WnR70efD
ng2wT8l+pT99rmgphdjVvpruGfgNm5HCyaorNFXqZvHGc5QyBEjLmxtpEUM0ADgv/JvmSyXtdadz
6ol+eKKbPPnXFpv8HWMRkLdUxDY0dqfJbdggu0J5ZpfcKnoX4ek52XtqDm60qvc98HJdFp2xUh9v
Sy/Nux+MvKvFDVpIA8cEoV+LXNLYX/Q7B4jzNWum6VYzPLnSCy8GIbEpnDDjUCBID1UumJ3a0juE
FrVBNvlSOvHxM8lFOmYPoVl5vvW9Lpnoe+0n4m0lzO3wK/mbrPrPS1a/GEyQDZfpKT6T3QMZ/U0Z
bh+LbsBECCKXpXADEiKJg9ayTv4qOY6fpZMb2fqjk7AP1isv0fI1IlVoqarJCo4UWOOy5PvqWdAd
VbuQtM418xXucX87lBQs50OUOgij4TjE1pcFiYpuZiMU+uwwQ/++IyC5O8MX/LyhIwYmkV6v3hjJ
2olud+rQWW6Wl2Hy79RwExb3XUVeww9lrWPq632lzdE8s+OL7f2uAGmeP1jydvtaQwHi71mzycT9
KCM2/xhXvdo7xUh8Knl9TPUvn+0DBc0oj6ZGAwnsIv3m8ocPRy9tU7PBP4IXUZtUAbGVRTei8F5O
IvS1cLqqkpcArYsffCJd8q72uSLuYXRqCPvWC3wpTNAkrTrnoWKdaXGMt7gims6bhwjjy35RICV6
lCicWYToFsHEA3U3W0f0kPK+CGHIWl6VP090rJm8xinQFxUa5D5FjklSwfXFt+NkMe+REJT1fVkV
ptLTZB6GNxD8i8TL3U7bnpT8DL0RJhrzE9D30+wwAMfqSK8zWgOOP5X6ZCw4LC+OS2eC4FYoHzMk
9qHjc0X1DwSh6oCPcKlEtc8CNwpFHC70SL06MXsAWCjxfrj/HfhTV7jTOOVuORRvZzKmW9leBwcp
yvchAXoong6HZBI82ESPNZUZDB/j2kD4M6STBToiRJMlTSt6qPFSNww5ps9vfqJ8jClmTXLAoqq6
4NyZUyqae/jTJHYqIAMJXWHeP3wyUATi7Zj1dgZROjdUcxJ+Hyv8DcAHvsmJ4qnPCdW1ZjUSAj7k
Ntn1ep955RAw2IvgnTPyKUwGVdT/yRrYoYYt1c/QpovDXiZDx7X7CVEEc3Hc5NhBONYZyx976qOz
q5ihoGQ/4rhrOVrncZ7O9/bTpb4f/0x58iqkUsVhXVkK8d0lTkwakkNfynot3vD5iaoYn1mAS3T8
0T3mgQD2AlVzBtF5uCBfuncG+X+wxAlIcP2ZrU0m1mztUHdWJMHc13hdmXhgsdw+wGFTDhjv5AM6
r8ekkN1FS3d2+n2jW60H1K46RZVxd4N2w6zBEkapqciDAUAPzmN2ivaGDvgzFJ4M0dEkxwmPbR7N
X+20F5X9vDYfUFdkSwdp1G3QmMhmj+SgKQjyyJKXjmLQq5UDXlyxY3jYWYaqJ1hlQNVN3nMYK0k1
7N3CqvC042V8XD4tYmnAnwRaUvw1YqnrB5rK5Q+rDIqie6noYblZLuAJDo+L+XuGlsjDcUdErGw0
G757u7YDuOU/QvSgyGHfQsHykNhIq2SznzXwAQgVZm5l8SSH9QMOGBPb4FpzEpU8jhU9oFev08TM
C3NDUO+UZQKuA36VXRv/evRzaXQFO72IA28y/AfAO7Fl+01d9IFNA8a57qVlC54SJT1j9j4VmjlH
1jaWllVivYbizTZoZdMC4zlBVUlYpxwa8mtimj9xXyVueeOnryx1QN3QMBVJtonnWzBAk3lSW+jl
jAO+tMXultJ60JsZpHs0gfJ2cZKOAt7wa/yarmVGyLO/2nB7Nbte9ITvTnH1TdjMj7dIBZzIG9Ny
P7SjoQ98zIZqCnkx74FRpR91Kctk+iwVKGcZw0UFm8TT7W4KrbOUBhijqRK06MMyTYxTjLVoFKn+
oxYmm2Q4Orzynj+Ph6T1GCrkzYc+cgdfV5bEaNYyUzZ9iODDPJ8RJ0N5cr0YHeiY8tmPtiAs084f
4f+qr7A2FHgk6X2bjSuPsdt2AbLQEoz0k1i8jed1UGx75PXCyBHSI/s8EzEsOiRNPNvXOkPhEVZb
0+kSST54CHw5NjwyEVkELEpEsDBkJU1oMs58EbNT18qR5yQycgSrM4mVLUpSLxuMuQMjvQ1YjULE
374vyvhEhuOgaLzjrzsgXvqd5FXaDTGrg3NnyKFeIUwsHuM1lUuRZvRP67Aw5XmivN2Z7umtXaiB
iVd8rfl9QntmvutDV4qEAtjGERAlqdrE5JNUmJcN7zMUYtkBSn+jsddhsDqCdb1Dkue8eV7FEVBN
W3NZnwF9UycIYhCISjfI1kWfDrrO3AJvcSF6dA0A74IDbBgUCBegTNj9E4ybpqEUO1pxuzxSyprr
QRsyeKb4SWC8YlkJ7GKgpRpsvUes5VtaBpWLifqT/drpt7R94jaGonSykkFEwJU9hSNrXP9iPC0B
NEfXt6j/OCJFNCBNRpjBgWjKBGbeECW1qMc5y3JkLPPdRmW3Lzh3M5jhwe2BCd4nTFxNeDW7tQFh
MUD5fI74CD0ETgH5E8nTuIZZMkfu4c/ZvtNajvT4zRKECeMT6qm01jKMWb1WI00tZ+nfsm7lHUJ4
nQnDbBHy3Z0cMVb96SXyjS1V9nCocI6XHNSGJpSBWcZ1YbRLfyRsHQsHzi+CQbU3Sz7fCPPSLjWg
AgOPN+4987z0JGd4dmBejPNjWP9uz17qkXrWUL4702ZvmSmnH3Q1FwHxvu+jy1L5BfEeGOMwCgHk
verClXyKvY0FoHVdVOWkbydXhg4CsT3FxJEB7+BSePJ9s4HpNHUPpQaujIc1PpLvF9F4+UEGW4tN
N/T5l5sMIbzbb0Mw6LiIHN/LGn0BbUv5bA/O4cuOuNlW4vwj23sVm3wxbehTHpYQNyFFuOMrG9mp
QDwd77+w7kuVeal3MKpIIutnSimBTMOma5uIzcCfLtHWOUt7zok5pymqvvSABU324Kg6emEoME4n
4SQ/mRjTOw3eGqfRok2tTzu+EGJM/He6KYDyiAsk1noHilrzuvKSCWAgX0ZGSnSQ2Off/selMnFN
u+wHiJpU2rSEAR7AvNYtUB6WgApsFhgQUr9zqvUtjgv9ePwEBYc4zDA0pHH8ZJGyNyU0sh31EzZg
ErhXWU5ZU23DFtURuy5PfFMDDl/MefL3/tvgwEk2xvpQIhvmv2HykiuFK1VixyH8vciwu0VZfxos
VMsEmQRjwXoaXdWQC3RafQ1zLh/1nDG9/XdrJtZjFNGJLfFyJ7aA85gn4BonXiadMWTHyRSs7xmS
JQ64uSU23jETKnx8r7+25NBNvUAcvL3cdfvRckk8sMa4MRdoZ6qIfwf1O2OfxGm3/8QIQxSjJa2Y
BfRP9bE75dQ+eKMryV19irvitKfj+Smb84kRliNQdRXTfy1VS80WOTDobPwYVbjFD8DfQGW1Sh8B
jh8Afv7OMH9rCCzhTFwuqE9gE35+Q/dQwYp6OFmi4KnVamimuWJ2Yegr5vM5PnQYw/pW/cUFpTKa
tKGkl523DVPA66V9rJAYKPgAfHOa7MV/X4W2QJO+yKrlApCWX3ORmXo613roT0d112KEei/FwXLS
ALyWsT9VuSkggk8mhobr3SXuy1qc/nZB6AlBuLG3oLPO6FbMDPY6ylj9FXCQWhOI6Hu5CegJ5CZp
7G4m2Fa1jccrm0MP/enZzfkGMzKrSNU9OmicJb3+9wVuJdkGUnu/q5TMw9/rGsksRdHVyPYMeWZR
HbJKBBnD9w3Irpk+EZ0Chb4CUltPwW8lIQsDrldX9nYY2JBK++RsnVCEJPHMp2QDZVD0NW7IaOuV
xIEw4NnxHXHW+NIyZ/VJYNSoBQGsxeB2AcA5eUxEwjILyf4FFRkHbCe2KKVcNggjCAN/57qbnwqo
sZsE/ANJxo2qU7Fz2HYavMP+OD6EcVHliKukGDUOdRibytxiWDRS3p13nQp1AiZodiyqzEydqgnt
t2XcQ835TuOCEP+7Shj02HjxhDhl1shDT9D5YYFfpJEcBo/xQaQa060yW0RdguaZmzfb5wnxBWlG
tc3Iif2uIBbPmT8TkrPrJypogRw0IeFRaDb58HC304X4DtNGmAUG1PBt8hVpy68IT/1zFaF8qz9D
cjFLB3y5A3mHoxHlYG0o7tlpfHg6cdNokILeY0zS5f1fZkttn/i/JW90CJFwV4pZacoWwUaNDdlZ
S3L89BtbIIc6fFZCXjXXLhG7/RRZTkOA8gVhx6OU6XoCy86WhihOVK/y1b36wsblNtvh6EUyZQXg
yBXWG52f3uxysARgqZNMoyXa5N5yVPxFDXQVDIAwdbpUo3dUqjKOHkYDVcpgmfOK8Sj/tDyhI/sT
ldx9KG2A5kusEE8moMAARhxA8z5OP5Hg4NIgAHjnmNHQMAdnpHfAszgJa8oVTpu3AgBnowSJu/P0
iSXFKqtf9EfufqKyQdUDCJnvqRs4d962LfoZ3C6PUDgKTWtvXhCkgq4MCodUdrHXr4kUj1/Dm7mN
HcvZ3IbM2lRqtufw/ci6yIfuDJtKhIwmh6S981z7OT99XynWYrHaU+IMKPlz5plejHrCdAG7QWWb
+WG5vGO3plg6/1ifyeFk50HgsL2E7vbnj6DR5DkKRxuxWTVcJhPgdOwrdnJC3LB/Z5Dy5QhAorR3
GbPehvim5qvV7xK5j3q5xMl29vQb+Axir5zdOqXENLmrP3YDUfgZGsO7xygPbaVKUzWNZlr1/A6U
gJ6yNjNTiWYrOaNEjfYUFCnXYHIVak/056NVAkbnA4/K97T7V3rdhs0am7VThR1BWZuAn48LY5SD
27pnCCVNeOcxhv+v3UzjjJiGbFCkqGtdCfy6UlWLaY9Nc/w7pevWmqlr5IW2bCf0wbIH1IsSYoWh
ktxeEFnAtc61eh8gFaMiiOYyjq4znexnlkTbQZmKez+UyJcLHGDro/EXXKPkn8JlKvD9zczXIrUs
wiP+hli6zcDb9NU/7FsDu7obq9tt9cHXVZMCSf0O8oQ35o4zF4FAOW7e6jTNjpkcA6WGhH1i3zHV
Mh9avBgC1ATyw9eVCvmiOTD3SEKup1YRMF2vCgh7DoxnVfPxeZXe8d6ni6ZuMxg9qFBvWFxn7T2e
VWh6vvQV2HpG86Py/G6UvoymyL29JvGy7EdQ2f6WfszXds1O7ycpdEAr6J6vmQpESULWpLEswd/3
1jvED7aaKtzmfuuWb4WVDagi31JuETuPta3Gzt6tMlEREZ4r3ea7uiZb0kZKwLqgsUz7nLBTr14U
jjf/s9AngQQDO38/WqrjACj6zQOMigHySQU2IGfy1ayTRq47BnkmvgxlWNIPBaUVeiGiIa/G9r8e
nN56cmQBcdVee3utxbZgQxnQf+r2DvYMiWcY/J4FkFrGYCiBvxmgCoZcwSk6OkL4BbW8r/kk+xsa
A7FVM+3G2lnsIE6Q/rEH7GtaP2FBkyHf5LUzyM+yuIY7DEWqyECf/n/8xv8Fl25+DwxqfaEz0KQK
SPUecJ6slW4RNP6geBgu1mnVDMbQl8Lab+K7wBQXJWnlbYUqJdnCt1U3orU1FKIUgEs+n3Y4Xc55
T7Xd41mLTS/nN0OajMlWPAUhqXmcX1+PuxjcRs4/ldpfLZXx+BV9KvkpTSaONEA2YtkoQain6OpT
Wi7Eq7B08HmMWuyMbe6VCvdVUFMEkSnEf3xv11BBnlx98wnmOKakmWu4RePWifHAXamEOag9kvgP
3KcXW0YG2LhJgNtMG0TwLK3JLgALrXFcgQ+L0pFjFtZ6+/3kkYmG/BT6kh6XO/zMzNtpNlCLqO3E
g9XO90SHGZas2QxmsY0db4dM211IA1WRvn78jNxvg+2dL4IjwlR23QR6cbQ9YRmoxwoWL06t2PkI
O2goqFTWAdlRFj/SPSj1keE+mMKm0ekMqHV1uE1Yqti80t4mhqdJtzw6jIlGJtBLHFKkWFREQE91
+998l8UnvyxmGJCFWMfLF1J+vR8IM7f8z4/wo5HBrTkxVzpEBOqZXT5iFQNIbd272BuL9/IJwgKz
hEjz4a5497pC5Kuk7Kc+WPdyLtF52kv6BCoKlUpzs21tsL8Z6ASjKhTNpGNWirNNNXAPvZCxPR+k
iU+UGhPWH5tRe9g2UfuZRVsQVL8uqacUilci/pekNOgpUEmgGPEcXxxwOPUnGam68QpuvZjHmRhX
HxgGdbtFcTEKqVGe7zR+NrZnBQYa8/BgMrMAwvfmx5WpttyhlZXtCh2TIqiLXTiM46ibFatGQJiX
26gHtBKAvclJHbw52nM2gJAGvyZr1EyEmYvaw/ijbUDH1LSZcSVsq9H19C+V7qWceR85c1GaXJce
Lcl1s+MoXolLuCDUUL4HNSn3kLYVh9UPAifGWSFEu5K+cIuipqtpd6Q7Uhxx8yjrf+LvobSCcrpw
oD8Ianc9/9kfSlKQ+fGm4cUVZQ0UXuYc57wkftXn99SOlo1xWaKs1Vl+SFtxk6tcPi3oWeC6lXM/
qvzjLcPEBdI7kmS/V4Ixp/0rTZ73hlcD1WN/purmDPkUrMzxVPogPk5hNCnVb4QhwZ7ZarLexLdN
zcrsxgFDVklmU6VD29jRh377FiAvZjXLyZJaY8hnXGbDnzuJ1v3tN5YF3U3u7oAAiMfjgp1KChsD
5dD6MEf91uVBVtnkJBpQm1oeDtyFlLfs7rCs+7OmhIhWnRynvvxo+RA7sLlCLQTjAhhd2gmQFolJ
XaL73fNZtRK45d366meFVRGF58BP1J/AYf1vVT7AdEydiWQhSG7YaWUlWNtuXOFvsKv5AKBF5bD/
shFScJCVqGAtJnmOK//Go3OCNiFcK0Lom2qYl4lPmJt1ER6gkJkf4y8U1mCa4ainkLxumEtcW7ov
Ymr2e2NBlfutCqZrNvW/phPJBOfVBJMCmE2O4rd5LdrOAsVMeVHeeA342GRbDvIu2/ZughS1RMlU
OYADivrRrquW2iiVbR+cPwasPQdGcAf6mq5J9aWkylreOld6J3uXAmyO6yI1dHAo1P8J1+FaT4Ob
hPHw98rb4LRmKZ7RAVAyz5fxM2rZx25wdjBVKta8izVVEbTw5X62298sigKGFNkLE7DSpocGkEh2
/XT12Or/73lQx42jccu/pDaTWHQehFq+0fYFjQI9Tjfuo+aaqZHitI2gAr8GlZK0z25TIHncnCl5
o2DqqasRyXbg6vAH5rrrqJvFd4KOdFEP5/Tk88l3yegTAn7zaJhiTOdY1Qss+aTC4FwWE+ZcRHy0
OpmzCO2dmYNxIruz9iYFrXTNKUkFnsEDKi0IociTcDyjpUrPSNdnqaNDGRsx96+wl77bJ5Hx0KYI
PZ7koWB6Zg2YS77eKFMD+2gMRwgixvr+iNZ9AqhWgJBSX9MMnqIyl6pAZ/G7dFrl09ltjL7a6Sjk
5ES5DuH9nAHjARKHKEOgwqKqHpuq8fTvzhcAJlg5ViM/sR/c3d3/Q6/ayHQ8Vc8SjV7kTmUZtYDY
NZ/SrY9dzXjAjC2Ot4rCRyZyUKJKXxQWup/qsuA99mtMVqeu3v2kxaurI1RfFF/Ade8LbXEzjzvZ
F0kfpU31qpQemFUL+Y3hMv7dQsvZvad9jjNeED+SAx8o7w0lF+QbDW9BnFG/q7G301xIdIgN/NoA
Jom82c/GOMzxP1NSEUg9n/xx3S7g/8/VE90nf/uVH++4HJHV4wvfdGwL85HBloPaZ5jnKvA9f2aA
anIT0JogNq41yHYspFpYnClNASmLvD8ORCHD+pxyslCHhOmFSMLBO6UpnaNVh5zXXDdLvToyJSQ1
fozemJ9CjlUDH2yLQJMW9uoEPptrkDjIurmEBNWahF+WdXFdlEA4eqBnX4Bvtmn4mB42b+ioEhkN
8Yz0zvzqET/yWbvvN9hKbzOoWXCppwqPNhfv/h4/DAo5EWaipwbgMYU98YLOvHCKSlL/eR/qjzkN
ntHc+5l3kKFMR8RqzE5IubpdutH0lkK81kIMBefmRNA07h/qaoZm2KWR9Kt9CQzewZHiiryY//x+
7JN6syIFFcDoBkmfnuMEdpsAoSaqCIgvnNniphYfAusruCkNYPR+P0OeS8GGmN75Omllp1muU+oH
470MVvOAhbBwMoSD1Yfi3dcnlmRQGvvOx4T5Klps4YExQ77C7I6l9SXeJDysieYGPj3iIYD9gPnB
Nx33IZP0Su46sAhgCoe0TiFaJ6MWrV6jIO8q/yOcETl9zIiknJ4P3RWIkR74hVNqfB8t0U4ZjCR3
sv6lMlR5PF2nY7i50fwfPdoUw5UMFoxqLsKvvqW09+WLbxDQRe+lDbj18WRwjW78LVS43Wmb+s5h
PfWRAXYs+IahsQAwOV/3EBzHe6/UtBenMJJk6t/uRUeqZOrtek2RQx+SELc0s3NlRTfk5J+E9w5x
IHuGufVXqDCpTy/rQbkFKp07QgmWZ/UG1lcW8EBT6MVKd0p1f45v9StZ+gvtGDqL9TcpmmiVUFFF
V2DbTB3CigDwYumbsvisN1YqKiebrLxsBhZzqfh94xSOg3jEN/ZdAD/OY7jhm3oMePgySrILv+U8
1idMb0JQMUVFvpBthX/NZydlPArnTaMZ4DjwtjXJd0VwsBp9vUpxTpgfrRqalmHBZZiiALRNFMpC
AKOIV6qWkfBXy5ynKIeyB5dxIfhckgMDcEA/jUFB2s8ZszMAtcevCX5Nqq+FbTwoc2aUF6hIOmvq
5ah4zKzaN8044+vD2/BU03umL8MoLZt/ZKtVojJPhVPEQBvritGF9Ly0iHAjjwRpQH1zS3WXaL+m
p3o09feTY9l8DVHkJePmKZMruEhrNyIbxthmtwitN3K4oC3WIC1qZ4B2qyIxguQAEge2EmGcSFX0
eGUUwhMqsnkTZ9WRrfkcS62DShrdGUKCCsJZsph4f6MtpiG9K5fUtD38hKn5perzXbcM91zckq1p
2ZGKApKsnGi+CTfVtLUJzciLm+Mtsk9c+8ck27BCLX/ts97BDcchEDcGWPi74J6CGEqtoyEhTyEl
UA/McVHjRHvlp2szZgppogHGyBpbQIgizD7eM3y9DNn1WhbqFVXHEVaaOilgfLrGLSqatXqncu41
SEWcAd41wMKpboTSNQITvmVD6E0sFS6Y7c9+aVEnIkW2G09HGcy7R5XucSOYfF3mIMI8jHEDJmAD
ce0czrgfsGrZtVfUe3fE4YG4H2bWHWIHRObAC1KHoDTdeU35sNP7NFjCMYe8Y7Jx0Jy6OaD5+MeM
A93oOfcvk9voGn3VpJuM8oGXGnpErzcwEI4bJPfDpmkhG9cVVhyiaYw63FyFm/5BFuhXePSwjZn2
Dx7o67EAPND/fKMB614NLhoKcy/HhGXiEUiZMpNi/YfZi+e3jCcA5aoUy7znM8t7+yxSnUztahqY
GKgkTvLbI6JrXtgFK6x//kY2skJCH4W7E0KWw1LyRUlsY6Dm7a9eL+dEyeoCyOfDHPX4l87efu0M
dgLLOEJgYrI6Tz10ZQFMAgZj5guX18BL/K4kM/ku75zifwGZx/7jcYRUK8morO2Z+LLU65uOiW7Q
2UOXketohDyiVvfPCQ7auR/4Zg4vgEG9LcWCx5nCmRBd0wpJQ7Bo+NEfX2UbmQeeYyR5msLW5taG
MDmFl2ktfWHrBbqdy9dyvfQu1fQiZohcxESXbgkqKMFmeEp1Fnk1Au7B4WfhPkv9b8ogKYvuQ2Gu
48kb+KQ1yuooIa6QPrD/VdE4Rd+gjQwR5x+H4/hR/qqFijSXUD0Pje8N3W4clpjD4+1KlL3IYG98
w/rq1sibnE5r7OzGnBo05Z6ePUmEfCwtogGCqCXnN/pmAVqgeqt3nEK6o1j00itEeu09XppbXeD8
XwKpL+Z2Vf8kV2u240bud5y8NlwmKKaFsjp0MASsG1g79oWqDrLoZhpTKpYT9KC1/mNXFdj/qqf8
6e6XndjcouVLzkX8F+aI23V4spnvBxquKHQfN4574cLCatG3vuY52AAeewzcWzlBZFeUlDerzVlq
fn+4R81V1DxUAGNN3Cfdu8HHgZq2z1Ie9f+RCmUm0Ya/TlWqOOA+dnUR/P85Ab5pkT0owPOCQaXI
Ht54kVjSCKaTJpsg2527mZioiQsvrnxmVD1ICQLrecoBRHGadIBGpQzivDOO+0+8PfoCZM6L+wvI
KCcvJ1YJS9J3iAAAqMN8MnJwKyV415uqAdlRH+fqVxerBJ4KE+cJgli1cymxvJfuE2xiAjVDHJil
KelvSr33SpUYmUhtHdI24CVq+6pbwD5giLf/ep9rH7Y4J2G6XmVma33a6c4NugpScf/tupdikYre
HhabWaiSie9H2wOCHcKyTpdspWNIuFQFtkjA0U2lnDCg4O6LanQZ+7YKZ76XQAjMhZgwVDhs7GHw
9JjN2BjyMBEALJIami8SsDSMBTwPFYdq5R1ra8FHEIQmV35LKi2oW82+sL+CFwKFOdDzOau1yZVC
76qtk+Khb/uQt74h2Dvqjk9iC79fDj/VNKG6DBTrVW6VNNW+uzNS3E6m3n+OQtoedjycUtg+VAkD
G/kEG0ygaIm5dyHnjQsLEiitooqw4q6RQnl3hpLHEL4yKB4zRyIEQFlAcdy5Pt6HRKK/OD1v4NC8
5BjeeXVxJpkHOR23JdFaRc+NbCXDWE4Wa/JNDaRlYgQJLQbczWr7BPuSmnzSPPcVBWZ7wrcQX4Qm
tGugNLtjlpTRsNWzwVaur5R1AJYsz0aoEitma1h6I78APFo4JBL0zM9N2T3R8zKmABF0GcFQBbt1
PJ3whPOdpxty0Klw0Jig61+nVHaQfZu1GI62jOarQZ/KzQ0Pnt5Hn3Z1ZteB8wVwor0O3DbcRY7B
YrI+zAdNFuI0oW7eRtTZOE50iItlR3TcoaAUGFx1W9ENz6dyE8qVctw+sO6i+VKZeKzsoB2EhCIP
qW3yWhVGoJakWYwvBQDNPjrNVNaGe9GcZtofJqV26OLgc2xmy3Z79IT4MDXZ7LxJ+Jh3thM+ZHl4
bGUhbYPzjfhwYB3snVhcZvkvABnenpOewSEnD9r66IVwA2FT84lQORXAZbIVVDBMIfCSBojXchg8
1/v1bNUdQpmT0rYCMBl6PSB1pANg2wTPqv7+qdMkyBcegvLZaD98GJvcs8k7PCpm8g3zwVOxnpsV
YBd6EA18nVXjhOpTrkJ90YELmImTSbBoBXPxyoSXvORNN2yoHSobBLdjXgnfQDXiqkG8X1Hk4guk
z595zE8kwQHoBg1jGKfZjMv4KI60hGpMshRetduaDfeqcOl+/QVEzMjlzfyI0+LdJihh0YoHLyOg
rXDg12BhSRC3Y6Sr/AWu+MMOY1cRxkFj+WhqaQ5c2LTc6HF7go0syWnDWitiN/KUYeoAyuBY22+O
4wFtpFhSB62DLQirfCa1JZoZK/eqPasan0nJfco/PVAcWILwme95VLZTKCPYBLUeBxrNKBeS8MBB
qIuTVqXvF+qDZHAcmmVv9nZLz8lBR6odYjnSnd6Wnm4TKX43ACdU3u/wVBOY635ZNvZ6K2ZdQT3N
OH2YFU6JiaOiygAUGBb+AcamL2RcN9kF7zbMHsHIXUWDv+4X1lZHWr+r0V3LzFr+XMqgn1zKH3Ax
htdkbk85bqRc8l1zi30wO9Qwa9pvb2Ra45mJdyEfMkj4zX3gkliJO2rxBRo+6rXdPeeKe+56TqWX
rXSKBpMIq1Iluz4KQa1yHrT/YRpDHkIuCxvY82pTERc3BJQSqifYdhP/JeaO9uZGt/V5NCj9+x1B
sHw1zElTtm1SbNdQ07/4BtgHnO6VceWrYQY9hWcl0Pu7pAcxkG2KRsXxGSZ3JwGk4Ev1Wk3nJVCG
wrNPd2l0l15tcLe5/0jbCIzOqeL4YcfOU41bSgfmFk5u+YkHcXE2blUdpfViSr7Ryes/x/uUgDYZ
8ohoZ92/c6PjNLTuT5BJnWh6o13PHkUajI7cnD5c8kPTqjQEWTnUhoJYZ0niHhK/PGrG6HIfDSg4
+QlBIhwexxSlo/Pabf0pDV2mxwbNJds8pZbeqtuB1KiISvegW8qwKi9v2FKrHD0shcRNjGn+zVVp
W/c5eTHocZpCVjy2N3HmiE6eC2dg9CMahlcdiPkrJYu1TZWpl5opCTIZyPHD7Ffg82h2hmt0Mjph
nQ5/SXQIrknJwGsIfY7WxD6SgMAnzdxMvk0F+cFEglXNlkAvtPtpJTH7FLa4BYJ8rMoejp/NoqC4
VFGUbKvi0Qf3ytvKZoMHbhpFZktCyLTsHFdJv30jI2zG5GdxvLqDtp9W09zZFJN3Rs8bbhDPy11U
e6yhAtH+leU24TkUOpBYnFa+jBgKX8c9sq3+HFwlMlY4zmTTdNxRQLKT+C4Q4BQJFy9PgpzibLCn
cMm4Yn/jAeTLnNHqTh8Ev1Bi1qoToK/RLPkhwGD4OzKAyOC+VBV6iyVBh+2pcLlhxdcBRB0fr5Hx
C8hO8opC9IaiPO9DVsJcIpmT9UFuZXxWx9eXNhNH0qY9Q7raT8NGxGbn91O1kBf4gACaEAFM6YWU
iSvualDS99TaeVIquDhL4nGabnqy/of3bOZqD35XOoSrDPrFBLBvudQHMtLwH9Dgm/u8G54eioSN
7k+krm3kMgpeuD3EZALEYV7V5Crp9FShSiL1dz9qcCplFgV3fIsnScje27hMhzX+uqAVIx1MFhpj
xdZEkalqnoqUn6osfzDB36VCmEKt7mBq521aU3ICaRc1U+MX+LvI0Eg9KpmGiPUrmKwZ/4n+uAiQ
KHu1akDdzM0dF9x5CjAfFZsSbXDfRLBs2HTbNxuk7vQNuP1k2a/rP6PUxMKo601zIoXrbIMbfCPI
3VLRYAJrzS5K2P6ovuSfTkRarW1Q1qwH9YF4rFxyoMo4yOgPPDc+a80UcXrLKpRDFtLSePQ054me
uVSxpEC/rSRrZTn16VDHmVGYtLAMwCZeFn6WFiiGrJp1m9N8fQlkwL1vAE59OiKshyegO8srYvVb
FYGNVM5q5OXui24D9Pq6uNgztHHrfUkUgpbd8a8Mx8E3jyOxV2SSraNaApZWfVU3cxcbsvfVdQ+u
Q+soXOuf3jXAaYyPq69tY0r3dWxDHrJ6OaMcVPrPOiDWh5Qvc0AgyjSBFKtY4dPMsD7eOdhm8Fk4
Zl9LrEeV1KUURZ2MWDli2NVX9VcHSAonkQxVQ49B+Vy0IMiuFq2FvjXo19pk/9z4/Csto7QGd97P
B/5AJVhuHlTXv9quRlpKMkvIShE3dMnW+O5UNLkq0uIFQiy+z9Yru4zCVu/gDxXlrG+iULk20sPe
7EH/REyvDq3DNyISN902sOzSpaprK+xYOzm/P1or+gYSBaNu3+anIQXDXJaALvArLb5wN2R+ZfW/
0Br59hfUo9AT4ccycD4k0q0RnvZA9XLwNESyCifjVxw+fIOkpKh224kyPx1xG4olIpaRxV1iQTWX
Pe0wQdOekdjmGK1NlWYZkCfI6+RuRjxN5vIyPkGQxOwZMmJsfyAlswEYA41S8LgbYtSADQTN2dM6
GBX+rt2DAHUZAxkoQsL94f9o9di/nnhwLZc9S9gQs72ZZpc3wT7BP/o0NBd82iXyyu/jL+YqC8q1
aVG5DJk4UPHIUdPv4xLfeQPInSxIev6kDV70DRorcaasNTVMt54ixMnJk1FyGvug9ZJoNbgcVwnw
EovvUZxD4Mi8Epq5oUhctQ4gHN9qzCiLstUSinBPr2fW6JJEozM06JpJ4sj5lfqxhWI0n3qR7h8C
Pq7sbswqIjKoAakf1WlmiHhagKA4bUdQJyvSqKX0ayu4SLKVIsF4bhDhzSrXPwukpzKPSll6d7Px
ZwkkXWKprOusyQ73iz7395gxMOtQK8xEAGLwym8mVzWUC6qdOLsxLs46SjEjQ3Z8H/5+Nr/3EEXY
wfhIRs7FoaXIOiaO7g2T4p9x9YjhxC/FC6t+J6T7Qo8SToaNNIE5sgsq1I3d0t8SJ2R3F+15p597
DoDhx7DUJKmflbHpdCEWeCHQInex5NkrkE3Sz6u1I+vcaV4k2iGkBhK5dE2JwcPmSt+ejJ7HXIAr
XKmWSWGeaOHZL/h6H4QRl20hsocZrWan5Wju0NPftLWrStiikgbbPEeVJTxno3iM81PtcNxpmX23
qtVcIofucwkaVHYXIjOyZb1Ss4nM8dnlijbYvLOhXK6lFdKJG+gLk5mYegZov5o8qXqDZMBWzmgf
MNZIikC3pzls5VHwHBIGEAw0GabZG1XkEox8dv0gS5kKRNva62bx42CL6LjYjwRO2CplC6BLw08v
zywjVWXcd++xFUcQIvNdgOxdxHAaVC64hgk3uSdDtqauq/7XZlOhhnOMLhl5mF+rGyN1ALAyWhXs
qljK5qb9O495Ev2hhpxfW+zMNjftdTiX+ewHXCp4i+g/IXXAz4gaKwOTyT4bsTc7bmvVX+vM3Ao+
oV0bMkBTget/q/Iw4RH68EpV7jGgSqA4IUi5Ks8mmuHB8guvqregbsbJtL8l1ZGVK9zxqCYpyUYg
lnInrMLE1yFkZcxV8U4aaUtdcfh6FLTIMFpP7/41NDK5QVAYS8mN2OaZlrN0szJZpV88+y7AvVmH
IwB1Ffw+rZIAcJCuxWxSdXovFYf+ywBDICia5I2Yngk3Vt+acGXtk8GhEwp8H3MM+4XuVJY/0Ez+
+ueoHr00CknTBwUpHOT16bKv0P1EjIY3K0jIHz/+CU4U3LlJNidxULE6OfPpd5UHSRD+jXVp/zVA
lGTNdZypVfTnKXTf0Gtw2E4vDrZNkC77oUvbLOnvDlWI08Na3cZpam23wj3q7DVxbenB2hdJbCqx
IWWoo1cmBLmP5wur8IR9I6a47HeqDauwbZ2g1ov3vXPB+QUluBkq32VyhSAobgkLESOSea05/rx4
WSlMxI34BC+e9D5So204kkoPW2aQYQWNNh71DyogzgqE1TcFySxX20Qc3dLW3BUPgoFrMaRiKJX9
N9DRwMHtjdmvd0zQDkNeb0b5m1TcAPqM93NKq9h/rx13koYYuHNmWoFcGDI/QDf9qA8V8U4xz6KR
TzByTs/4GxzEOeFgHYY46eYGL2rS6ZP+aVzaJK8VMje0nVK4ALVic3LTzvhwt5AYFzgh3vqEiX02
2Tb9S9orB0j5pgWdr9IhimOBusPEpPNRpqTOYK+vUiwgdpoH4j9m2knJAUns0rJPReBUlw82yd4/
QN1+8MkoyAr2xRQh7FwoJh+gdp3FnnU9iaq42Jbn3m2qp7jDtzxWaXA/wfhoeyVMmYA1+aUBnD91
nnh3H5nYXtehTONtmvKbSA0Vp+sU5pKZXJQ6OcBhMuJE1hGkmjNbeNkY3e4CW9B5V0AKZQEJ8kO4
P20zBLplsD77RFRL8lVJxztipXj7T3Itl/e2M+AnmMFFkB3U1isk8Pecg+9IYC5oVJ6EOoN8BKrP
iYO1LLOMAZZsVphHCaOpgmF6FyCoebul9kLI7tLKJ3/JbltKXrz1kEqF9Q3G1vxTs4T2r3hVIWsX
BFRV/Z1ZM8AnyY8S6LSKFbpetGaSe5DU+vFitybkD0PocnnPjoFx20ycPXZdG7HU1+zbHsbtYnqw
UYSmMtToA5zGSDT+g6fOlQUxxqcCMNSOTWtJ2PbADJtzSE+jrhksl1RSG7QPzxGKsRlNeo64pZkn
FQHGMuU5w2iZ3c8UosxN8vlhiM0aBPuZ93f6h6N0fMiAd+xXEZab/pIHHa2gIlrgwGmakNEJymnG
da87BKZJjrMAmRKM3mdLnP4lhhzv8O6Q0zWwoDGg3ZlKaBpUHe4CqWqJu4mA3yxV1i9I3Oh9cCl3
nsY7go5ubZTT6L6YmCZqfQkC2N+NXHlt0uTjRG5UMbD5ouWMEUjCQD/1S6uhxZFu/Goh0pt3DXJi
g8H2aOh6GNS45Fd9/tsWlYvEfba4PQeJhZQeMJGdUPUjuQRssJf6wB4GrM3IB2w6+2Oup4ZIwvjl
lcpWrUJbSMZf6prOPAS9MI5gps2MJNs72NjPcTEfBZxl8n0w8rimHLttYlV5/PSu2wE/2NBp+fma
/Zeps4Rw4s6l/SFeg2r+hzzokiLIrJYejnF2oEST/dr5QOo/TByzJXctu+/o1JqEmzQpobKo3OS4
PRKMvng4KpkUYKGa7bNTr4joRxyCfCkTBJdFUZjRSpQ/gTmSk1kEBshwklf7h4IUTVZBs3OG0vD1
520rCdcuJCHlnh7hXOGfL0r6jhlBAxEQGPr55sZZghkWf03Vyi7Hs+DHzqLoogQDZmL1ZqptgDfr
P/xNWLkhtyuFaXxDGgcMGvBOWWMpRRmxGm0S620tk6vmueP5i1pPoA252KkuJGnSB0WF2jU97BVC
nLO39KVPyPO3cesE/VWGRvKJSAOHwze3Xp7oFaQ+R0chQqBZ/X+ebt3zJPF5Lov/8lLuh5R7oDfx
3lHSshVrmT0BrjJ0euZTzHEXiBmsQYfuKxQqWzxla9up2sQ9wLRVxO0vYCkkEkFpwrafSQ/jTJbq
1/sZxShh/ymIfuQ4XsTg4iLlPqFq1avGRiQCvrPIMVDarPA/1i7EpEcljUWbRuqRpd7Yv5P9XLYR
GnMacaX7Yf7/eS8Oo+kuQLwlDjRTJKGxigYE6RUupVQux/hPY91zeqzfKU/XcFO808Yf3JN0p/aP
NPk9oeLHDfp/U9vNqp9sTRVB7Nun0bHNddOFBEqtSOYKjgkFvL8bEA+sc6sdcvq2ERoJmSrw0BD6
lyFjwHPo8c29HtwQrXq5JcUgLI9JKpsQxwIqyL9aCLP3Ce4nfiCYW5FNOsa+NlmgMP26k0Zpo641
1Z1+rFgqPTXspW9HkB/vdRRxZQlgqqBZpy/XuGSg2wyeSwLDy+FexQ14hc6ah2F6oZOeakUKNmVy
hSfNbkivxo02NNvVebRO2J6ebpW7Mm4cqysU5dO/AC9veSQdmWafNMnHU7J9/TJK69GgR44l1pzh
I+1Lwe3heH5q9trhD6vxnQwpX+QvUUtGUq62my3z96fpaSGpUe9jYhnNYHv4OTH03DmRCKxLKIB+
KFVM+yhh1VdyzUdaGU7gjwAClChuY/DqNHl9bWZ7VvN8MpKOsbYIGySXWu1bQkU9bneEY7KH4QnK
xkdIf2mfin+doh4PWnvey/9Itruo3gUp6i9KnDXi+hdLJDxjcvs0erNlewzB0JgNFNj+8WrH9+dI
TqpyHz1eRfqSCXhPUZXa9iTa3vPOVao9W4gsvUvXXrfbN2pMGVFVXC7ZHM/FWx/rXScvHLmJN0uF
2CxALAiZDynHA4WSPfgosBpBFRHVsrAxlxIEa75VIjMpHeeAHma1IpGGIcR0FL5T3ebA1pjmnR72
CQlElkGiuTTLb48tB4KkhAwETDgAuW299MRI5THSiguLPb5LMK9HIyIwu1kAmGE2QCvj4mZdjQRf
8g/VPWs4iW6YcWeB3UMSAvdmKddbYCVZ9VjKd3ZyD8H9+mZenzhZoHaNiyrSgCv2Ku5ADaN2c5UQ
BDPXNxue9PmVpzUqyG987N/sdDmPDUqB4WdbmN5/cJRA3WRLUL9DrZnurE+xTSUt6KVbRQPiT4wu
ZSxn24XJjQcinCuyOWP6JkldgIioJpIGXZ3GrnHNee5/Do7PwIr8pqoun0OhueVUca3boJLgVXTg
Yi+g1JIphZbpPdQWPTeQ4LLu+64vuqiOv9iOCadhO4MnL/6JYrDa2EKkwvUGaXY0eDV8itvf3MKn
gmJSlVKAlxChfglrTdqp6o/T3JtBz4fs7HlkrczJMmM0JwLW1ndz3WwqlC4Asa1+E40uUN9AfwFM
tkODKpPN3XwfzplUcLJEDtWNsW++Ibea3MVcm8QfXCp13aiOVg0ba9FRQc3ZJmfuCJUITAbgJ3xq
Tc21z6jtrkwzFv1gNBkEijf3LG9Hf03NI6fBJuj9a96uessNzmx5fgB36OpyC/6G0p5dtvJU1n2d
zwpYP7ttatAxy/40bmPLJmMD5OHnF9eWQLm0IW0ig5Ly//qtQH+uXi0l6uzX7IxgPCjxm9PRnU+m
AMhNxFTHp2J7FjBocWo0iNsR2k16CA8ctwcR0Qc3Z9NZQkuNb9exFh4InwDaFewWHBX/mxRkTpD0
pJV9xgBZJaemYEs5bNV+bVfhNZjZS9euusX/LlGLaHrbDUzsk0MFPqVR/aW1SgtIOM2Zz2fv+0Go
NpInwhaHrT/jsC6MRvqqpRWiuvRDi2MnD5mUX2bO0HHgXtnELQmOzQRSwH7hipKhe2e2iLvw+FDB
DXkjY4+avKLDba9iGqj9ut+JqSzTMBSnVa29x528Q0ADHK3XlaCuNv2ZrD0YrjIyecNeaSEQ7OQI
CYTcjIBjqIULyHSAltKESJLBUy04j+S4PSAE5gu7cOhFZ3lWE1LiOasfKRlawdQBsbCK4V5mzg7S
0xQtAhBsIfZZaq4Bs91Y/S9P0ow1GmU3Iu6zNcMr3aFUkMaDNNaiki9w86KJlfcBYSAwqY/ic7uJ
TxOYksDPU4xW3YLq3O+aNk/K7J27HAkLaKjANksOdDDtSaLX+g9ufYdBd43zKYx71L/N3lOJp1D2
8ysd2OhEJGpQ46UjopVWJSUZv0jIuwcGyyZoEE66rKeF5Dsw5pzqtrktSuNRnRwzvtdRfZyXAoW4
2ofzdQNiuAAyU6qWkcHXy1IHtz4SHG1VYhOfBbyYUX8Bw3rhwLs4nGTWKZJYCozwiOUL12SwIvA1
zQ1Y7SLbqWF3H4zt3M9fz52o6MDsBgBIT3XppILnSIiTCnft0+hnO0hl3LPUKeFPaUiTuUTWrhpN
XT3y/W7xqzG+BgEYGFlUF7N2os7cs0Odadn8lPhpdyeXlcZkaP2npmr2b1ph6gcLcAPWAkerFeyJ
qxH6F6RTaXF0PjXfaMzcEjDlEe8l/wwv4LWcokdIw+s0CZ804IMSFlqGuZTS7bNdAcCtDbr9wb7B
bvvnULH/O/OIKX9DPZbCWgBZSkyp0QR3bBVmtQN2ssGl7OwJAWAQoEtv8lqIhLZXmpe5Tfib5ZJ/
6OFN793HnOdCQ4uHT3IvozM09ZM/BnLvzi6rIiavvESU9M7JO7On1g/tVQPs1EWDVSzttgOmaall
wXzGUkVk6NQXr86+7+83vJJz3DQHff/idOn2PGpMyQkv93r+VZIUurL5qIWRW0rGXwZgoeiNfAly
9INa2r9FiMv689OjoF/McGar7jdVVXz7tdTKli4/cuqfmcY4qL4AERfdoXziQNuwQL3X0o3cRkB5
ccOoYWuX7+iLNWQNkgQAbBSM+onShPX1Ig1AesrU6HNo71ss+md9jzarG9mk3fiUnU1ZkTC4JJsp
2AjT620xk3cA3kHvtIGuwQDOCovdd5vvM4SffIP4rg57/Lo+/dXt8JTZxuK5UIFsSJp79RwvV93C
eH+XpcrWoZyZJiHkjhTShnE+uXVTzF3us7pdQiyqcLBqQxV+oW20OfdaFtJBj1M2y1dBDeYWJ/gF
yZj4tBPU7nkxHPFHm3ESSeWZRR446rTl2LU1OpVx3VH/nq2FXif9TRxi98gtzSrlIklUqcpzbxgZ
MdC3P9yjiLwtTDg4Hp4a945/YNj7qSwdAOGl4yxBWpLIPg0H2A28KXxKXT2BKKft/qRE5jhQ2rej
VHqITDGgCtVglaM/fmgCSAMKIfzuZ91B64qfcTHCd6weRKruHCxPtiXxGNLpm+VEGIG6ro5Q1pwe
/o4d+xk9Vm0UeEcDshcPWd1Q8TXg7VjQLgC+OXUAS9OWKlaM4ehljVixbsFj8dkQCqEN0TLvtDkK
E7SWJ3ZD3viC/Xa8/fPybsfEKUq49YrE4A2QEQVaG0GcYjVy+pNDL2ohJVf6whdiCezEz1nUKbNI
vk1caPXhWiUHx7BmruVcmSWtzAbpO0TFajWMEXidI8Z2XnlEPK3yiww3Vn+zXOjqIt0qt5avwph6
0In4TD0kkiFpwK/rUNTI/ep3F/GI6ZnrKgSjezz2PgXtmbHg8UmAlV1S7W7H2SojTUiuqY4osIwn
/xuAhF3Z6/xfVAPriKETvH5l432ydQG+Kpc1hmCx0nbC4DyOZSBcFiAEIb4P+dsScF4zHXmueayh
UdXi0FZMFNLbt5i/VS9aa41rt0XA+xCqcbx3wLrD1DNJmF+eAQPCaShm5GR+ovDMdA87dsLk0HEt
mRp4ViP/+kACkosr9Dbgs01I97tFTDS2ikX5/cj8lMqVj+ijRpupv+sN7Xe+T+z5pJPC9SvJW96g
z9hRStcjz0VBaVDiVXsL1cQurZBV4zoJWq1kjZnlTy1x6Mo1TrZfckfhHsa4Oz2SmLtONTByrUSL
21QQoiquVKWNp9eT0+CSJkO4U7P1tyOVyle1zJYBrPxGc/J1VSRjVt1oCFBXZmk8KBnPMD1g77mn
qag9AU/hKtZGZZ+nB11sfXn7JyOAJMmnGFhoNAIX4PaCJJ4Vz4ovHtQjCN1haJA5F6xGzsS8GT/9
UpsfHAhNzcSSLLLC9b/Azh31CNRxPIZfJ3vZsPpi1pcZmqIvqsvjlBuRd/Ll51AKtcGW36lyn5go
jKWQgafZXf09LTuZb1o0JoIFo+PZEmqbpIAJXcO5D4xboJeEcZ3SxRL/J3zgPcKgKrIIFSkfwOAt
aXenktYv/79naF2VA6GAzTOGahdGbD/PXgr3zCPyEFz/Zf2l49bTHHlNW81MVddjni4llLq45Ohs
dCEr76UIqRBzYZ4+yEX/HN0cXqvp9i4PAc0yPg9tSwsc44czHKs5Yz8TDqwS978uV2k2Wwx00BGr
RORilUdJ2zVqWe6RtEYrsfkwLwNyc7wbVXmOeAZ1h3ZP+QA7UDTiqq4yny+8f33tlqtFea7oWWBK
Jmi2xYW8ms1GjI4ZLjX5oVwWpZoEcrgoapQ5ie+BKqO/LTw0msQ0t9rKcO+QV427FFqkktCjHj3w
eoMZQw6D2JPnX2TKUSR/ZaBkrseMKkP/X1psLx2ZxKu51Klb96daBUh+kd4uplYAQ42xdSHZAGTJ
f7wckuFk8fl4PfiV/LbhErUNKgUL9AOecBisSlV/aCf8VZ1EahgNIP5+7hASpjL7NxeAcvUoMCRY
pJj6BiIkWSUbg+Bzf89BkP/rsV2XDT/vezBONB0bVLTx4koXCIFa0f76F1nybHxjzpuvjCL88ZzZ
CqIzjZmTcLTCwt9MOfgmcFvHLIcQ6phmD4TfUFHH7eOLOSKscOE+fyuaL5ZqZngkURZ0LPgFUY9f
2ei4nLXqEdECSkUu5vea2lYxr8Qog8ghQiGCUlbfUmsvbAOHE+gC81c4/EbJoHBgMGlwV8Hfwrmu
GER1cnpKdSwsPiErVcidGBKcr5U7H24lM09YgCHUAFYtxSAAiNMSmSWQJG2Y4rjVoDKY1SIb8hZq
jT04E4MTRuoptxGLIfsTvMN/e+iAAsRsMtrqnZSUARWNrBJq6Q5FEwl/e5Mfi8vwvQh7hoxAKglT
r1FNmNGEuWXA4XZkcb8f4RSpw+qGeZFWNWPvFxpOE3RvEtnQPF6M03OO2LlDfIhD9PZ5XN3x9n7f
JwGk69H/Jw1qrlXQKbPXiYT4RDNVa27NjCQIh06je6Dk08e2WpHGqN+UUETGgiURzLjWrB4SIuKf
gKeMwsmSJX2OMH/Cqj8VnRxGISjSHu13BxQ4JxtzWX14E0VrpA8Gsu2kza/00A821JTtQQI4LO63
DDSyJ+VApFghrMkv6Djlb4snzHtCJr+qOoCejRLB9c576NqtiVqEV3JTCQjYIbtYSE9hwTuyfBRS
VQhBuYZWLleJGsfmOuo5x7WVcfyinKMbtauxpKsCbjCFPE4hwA3Jc8bmItDuWo2gi6e5d291uZma
2vlhR908XHA2spFR/0SkbgcaH31hUEhO3ePqTGT2TUSAWankI5TIQdpQDIUf3iXQ4HVCjPO5unPb
bbK3c1uVcqRiv1yQrfgAcpx5Bv67k2EptmlihRCiTx6Kp2Pvcx1xpvYXTMuZ7YZcnDVxCyx4re+D
av3v9VRxR1HgShs/hxE/IV/Zy344BK/+TjtQKl31PJ9w+08ykLQAB7jsyqmU7YfwEO4O+F6m62jW
KkW0Kougo5PUjj56islXtscU4yQqUpUGFwIPXrhTERkbk5nyfI0GjhB9zsnnMs0S8bctcm8us/NO
mXOHwEkFBCReBx9FjOzP7/0zP/j3QL83fJ8HEpSokGuN38VVrQJafMuTj0Amxk46lt0fRm0INPZL
BCZXH5ax/TLYyHmNVhVq+OVYBRQuhZJ1XZNs1+kAj/Hkj20MqkaCRf4PYxEERm7vGw5Q6122EesK
mhTtcEjTrY95j7GadP4OWfWKF99jAlOijXM/oFZZxACogNRbPgF+wpMWJ1nGSRDJs4v39UlFY8y8
+co/w4VfCw7r4422ufclkM9NHWxifDZ04iEkyYvYuoSkSFuWdtBYNM4grdvzF3Moxp8zqgSmJYSK
qpg13cl2fsSDN1ppKzdxDFuc87gR0AvbmRt3NC5Vk9nF2JOkFZBeRlivv9gjTnT6YG+LxKAbKTJA
VHC4zMgzdfJIvH76cvuARpW+kgHXWLzMTq669yk7KDQ8NBPQHtWhIFd8ALDD7c5r/4lykA0NV+8g
IsikzLksCBHmqL6hfJN2QHseLzcR7nojE/4fktk7pmoBb8rmfwNtY1Cr6hNrlJmp0zA/mhg9J/XF
tatUueYXYDO39LB3/adgOxLiDreyomEfYSPjmGr94e0Rvx2k0kZhQEK5m6j312C15GSegXSZqXc6
j8JyX5P5IxX2iFMlTcadA1eXwBrZ/pX4bouxNtctn4EaFnWZ6NxcO0KAZDavc51rXZOVWcI2eaSH
lQmu3Uxin0484QF9nVaJPgBVTIS7T/83vx6JldryrAqWhbuHP+UPoVq/LWIRq+m6xWHM7lDJ5ti/
QRHOISQe8fhedejP8u2bTt/EIx8zpJrV1vLS5hNCiyVqTF4c0JMgNaEKv1McmBIBVaTqfIqLjoLx
gGU56yJVXcjsyesWD/gisvygOJSqKfcnN5LOfTRY/a03KDxON8biSzVO5hirDLso47OQig1WHnIO
iPHRJ9G1cQ3PpT4raFCFrnoAOaUS1L8u1cl/knd1O7CUsIv8uMuZDW1Gk+f2zXjI3Ap16ndix6lN
JTuItC4nPAHZuBua/WyWQSS6F19ZfMCqSCzMMVIggDS1To3+MZb1f6ruUQUgJPZIO0e6MQAvCbFj
F2VK/4aHQoJzw1w4cZNc9hAn3QaPGuBfJwVRy2UMXgCu2ASTe5aTHh5vXsLOGDDVxw150+6pBEcd
Xu+veMxieVHRdxf1HN2ZDWPHqZyq0K4QhW5/P+077x5fog0uVaAJzAS2VURhOYz+2ZXukGxmT62N
Ct00BZF8rP7g1gXmORNJrABM1xF03GYfD/C//JfXtVUMAZUMFd5mdV1ebBmial6YOgGYMrwNQ7P0
N2i7dIkoIv1azOLnKq10ckUDZE1t35DvLngC+RBkg7QI+AB1BvvEXWZfgXoynBjRtJ/ZimY+t0rb
LbgG6TQ2ocvd0/m+tAsNhIq/r5oBDuMmRkeqcwpKF5GjPhjUEReqdtEgOCdujoKYmGe65+KJHeP+
CSB1uBSH4cUQzUQwIE7mlkh2q4NkLayOGve/lx8/5U5Wf+ZZPojjrBDkDSfRwfmp3uzoIFcB7uwy
hF65qx1PWSCmgpxvcA5we2JwkTGqoTonYepAlckwDCGt7yss12fkX3PJxnucZVCc6LYemBf+cOqE
p+1t8j1I+YN0O78zdfNhWZY7lZlQvtmAjGi7xxpUfQp9rk4NBxnzVKdISRrjxQ2gMSfjMj6Vv1du
K17cpj4wjYzViNaGyOwIw6yQ5EOUU7nNjrC1PrOnAh5cK+zvThqCCuuFthg3vd41zg1lrVZ/aelR
uJEW5/dxmbOq0VpY94WnA82YD8SndFTWskgoed7myXanlOYl6nSKrEaPkHXNHZVNpkO/WBZvWxCB
yHaQmMjO+0j0YioW5AVFNCKot/MgCrAFIgtyMHkgJs9niLB84vQKGl9lfeL4vdhaGwFc29cganZg
eenrvBqnNeIizTbIKW+aElE8Ur+z2rSejqM6DFx7hLMfG4uj9L1AcaUd1/tpr0W6aq+r61Ti5Rm2
GrFqfXsB+1t5LFIIxTDQNBqu2QaE6yx9WphGIVgEBkUK3OA/H8Fpw9OL4qzf/vRFEEgwfes8AyL7
PMPJvaK2Ijx0pgC593clhoiekt5iifC+3Wt9iL7bLO2Dn5C7Ri7euz7+jY0ZkjZKYz9pIzPH2hZ5
zDnUETnpkVjtoh6TPaF8n/RPDGSNK2COjdS6bQAOil39svnEw2twZIVbJLQZaVE1woZuhW9/l2Li
ogGS6ks1WhbEv0gbfHnYqvWVR5tTqt5zllLCkkHNj04yQnc1CzPOkgfHZeDQi7lBFv6mSVTeOjjN
D+lRPtSJ4XA7UWUePLIDT40ziBm4E81iEJnkr6fy7ZYZ2GChjk1/aJAj7/+/s6IoTTxUXwgKJsw6
rML7imqKtABhK8dvtNzdGdTT2K5ur0MlpdcZP2JG+zQs3HEK+DfQgGtvpWt2YZWEDquWvrDHELpJ
6b8AxpFuKW3ZXoJKqjVZnHGNVIIMunxAOXfhGQmSdVCqIoOYVa9gADZQ+9Idt+XnTFt9OorFfOCl
/EBWWH35WJovRa+Bm41divUInFr+gBi4+0KfLZBkh9+zo/xDo6EVia4Cgp3bvzNZnPAv4RYY1hc2
r7gVKJAQs4RbRW1FHQLIprgS6ZEZWA43hJIKNp5h1w3In7cnRAkHpaS+GXHQlC0DJ5LcIbkmBI3D
ItQ8Fw36FNY1SOGT1ezcleKxhTksKeFonLzZPazVXI/r2wZTQUf66jmvzCOsHEvNt7EsH/nZCdIQ
EmfL1zMAQpPI0e07Bp0Sq+B3P4i5qOc+IPupG9aepHrskWYsC/TZYiwKFDOBtxhJtr43eoCShoU7
/+ztDXuxz48/JX/qVCNEYiiTp1hVCRpMCI8i5vC6YEw0Rs6Wx1AJyEzR298rreQfBCuReJi9HY+6
UYVWpQDnQftsa0z8pqx/Jx/CCtRtMM+P+jvUlBZ3fFQXD4dk403dzNlT1J5WayHaWMP4otHEDmYb
NMfg7p1Z1wBbpOkRDcOpnNdslBcRKgc+S5zjzIjuZ+11ojfQWrOLVd53HV9urLjY9Fz9MvzJm5L4
UxEJ128R3xN7XKnT1nv3U+SVjR8rrOcd9P1LE1qzSmPhxegD8wnzXGXazw9gWKvTIAAmo+pP8yip
RSlBJ7kuSYsq64Ra+Lxy1hKa/1WSUXoVJwEcAidaLwrg4S9Qj1kz1fW45a6n7lDPt/DbprFxmme5
GSLEk3ffE0UGLQqIdwbbj44SeDox2yY8jAsNl+wz2F7mQnzqSNQe2rDARreZy32MQgfjG550jwK3
CRWvQhR/W8ubwd17RK1+YByv02LpItOEWE+t3qmgB890KGHro6CVSS96ukrwnjUxdAEkFPlGCr3n
BllgRAR+y6ruy/9d1cmTgm5XpRZrwmluxIbO33FkOkHpc2xYotcU/4VP23lJ0+EWtsRJAZepYog1
ouVhDhSP6IrBYn3S35GTF6Uj/mNshx7BayhOkbaVoRFQfBDliB8ZV71pkL9aI1E2cWgNL9AkLpa/
LOafu6ZTJ28RMrueDj/AA7Ys9AGK89MWwknD9pzY6GkJJrNEPRXSzs2Qzn1UK/AZNKeie0qlh0NZ
9Rfmiry9SY6KOZLnGhVY+LVD50EKAR76yBIecmml6fwnTGHH6AM4gNeW7rkHTr3iHPbiOEYqJlzW
UTn9EraZc2Xc3AJORybldsb/N4sluPkJ5ywzlNGG4fETbxzRf0PS5JPn/4nJvt7rFvo7SQ1r4yPn
gRMP+eZaXK8f4m7NdNZ2bYBmDlwDoxhXZOyjxai88vYgPoCgTXKO5ayoMv/4UWfA7gzn0Hbb/rWV
LSn98uintMlqsLnMSPPRFbCzKf7fqpSgWSkfGubOt9OCC1qsWxKiC3MHBrHaR3fqaTYgDEPu/HAV
SrgoM032Sx11kjH+X+e2NqLYc2d+k17A8FkAepyrRWK8jblqvZcN579ifBEcK3jJCteMYDKbZRcj
IL26madKgvwKlnTMB6Gs4IMD+hT2cPcm3OvVk96sJCgoSSWQ8mw7UNNEnem5voNBen9dDcP4pLut
j9C9gM72MSvJiNRwoBYcuPHmNZsVETta/18Rabe0vjOfrM3Q7R9K8CFx5eHBI0r6rumXZMcpdbOx
MfBGMY4WqG2/Sczy9MtD0dk+8tsvgLyE8ZlYKrBUuLMIU6lH2FbUt5ffHE4QRBElXE66T9r4DdVv
r6+VHfcsJkHU+k58Ii/vsYe6qgFMCdLD3Zz1nVKLCx5teZWoEQWBhBpjoOlG3V+W6+ame1OwAoaH
3NEhUBCZaRpBeerkxKze2c2iD2Ef5tgCfm2pCEtzm4qjnI7hONS0cWYOn5KypLjN/IgmX3RZ0BZU
Px4mEwJ6A5fQ9hpblJ9jAYpE4ZfH8Y04bs5CX7RrlnE4dXSSASvYsgP+20iMJ/dFNvwZPAFBOjF5
/gR5PfFIhLHLb815DBTd8KeV4sAaUXk7zruKLgY3d0YH/v4p5fgcx6tOmoaEjU/Wt3iDYfn26xx+
tkNk9AFnxvIRhFUkfKGTedUjnPvgko0qKP9Et4Yum/9RYO8cweNpmMulHjuzavChB6CTK+33RM8y
MXewjTkqjZQ+vczbpL/6r0M91ijjnT7srQpf3lbzeKNFGh6fXL/f/WAdOkOaIb8wUlYehcZsG+Wf
uogjR3S112MAvkeqfqQ7VdC5OTO3t8CAHkXT0GkQlNE9bnbzFP2CiafmMXpFnDyh9cmZij7IWkh+
cE0zCd35FPf4Ac68oZLFjCulCbkjXIqd41UIvTpfq2adQBUfePbO7phz0Da8kDHtxi8tLMciAsjk
KtYyeEwdGlIFCK7/9MS1TNSV8lknKZb3lLLjAhSFR81CSdH1mvxoeDc8xL8GFARlVtN63rGIFYg7
CXxQAUDr3guR8Jjs8sWdWOGbMLiR3VXQFp50YVy6aDd8hVA0eSzItGN1bz4L/Hc/w7Zve05Fncxy
BOzupb43A8W9LhvZJrfLXbfBTAbUZ9ZwEPWzYxV7AUuYa1bg0Huxa1+DK4xgSNj2zfzyQEaxli4C
Yf/XNWw+ZMoOWWmeYdkjONV5u1uJf31GdFI8vDtX967Fo/Up6c2KSkAaI82uuS8lJdNAzrrjQiGV
sc5a2mwE2vs/8AheRIdkdsvQkkINgZPoL8onobj9+pk1iMVuH7axrWifvedAO/lGAiaEnDB9xeKH
BkNjQa/k04SLq1fBt+w69iECbmkN0m+uLslQesbVfthhA+BXKGyaGUaQ0Ef1uIm7mFpNuletuYSH
eJVEecpWmL5VXoodKoRhePmh5CJhanFAF3N66+JWZMNVw/FtuT5DrACA3AkHqKbF2AErvAp3fADP
eaGyjyiRme7rMN0nj+pgCPILmKqTU6QmiRBVC2OhAjmIf0UlICEOcSaFEiaAHsRFS1wCELEN3omE
wvtgeAlBC74Tu6MhlXZDUgFuLTjsUYkBP+0s81jk1qes1k7qzqrhP8z3sFpAvEofIDjErodIsPWn
wZCk+DTOj5sOdhpWcPGocieWkDS34LfeA8kNUB0E8eWxlfop1bfd6T+K0xOiHLcJJseVP9VkCe42
xsiG9jV6rLP5qE9rf9OCflFZE/A07pBPdR8oMCXCZkgbDBGs4B+3XoQoaIhqp26UZY381CTPqtFE
OoD7g1W4ETKKT460OxMe3ejQBl1Gu8EKlDdbt4Nx6EAt8+njUk0zI/VpmJ006xxPqGzTmy5N4dvR
fpMr0v5oKoh/OeUhmzU6jH3xA452ss73b+Vfeu7RJTSBxFclf1+c3qWQbt8ti5iJTVDu4H6jyKFy
2nErqByQ9ZphZlPaQZb8f0AF6i3UVvzy5p5RP30lNsC13hppqIslxi2wGBmDPH7KTnJGk7yzgRqI
ctzr6nZ/HcFBuAB48jGrVeVkoOULlA6P22UfQppRt9KwnpfevKe1JpK30uTyqBJwaNR4YPaGfFG2
5xK+uc4qBJoRZ+HZ6FbRi/zn7KabiB6EYgipe2JqVhV+Ub7V18az3SIcw1Zdvm+kgyqshzfRqUDs
VOEUPzDqO8SwKUEBtb10Tbn+EEc1ri+/pisQfJfVzirfD9Mgl2ePiKYxhWfPP5R6OA5c6HLg3k/7
oNr19upe+O9X6elkzATZ5VDiMJ99DGAMUQMslN99/AyzkK2F231PEtkL2DorRmHUX4M9Zm7yqsZ5
Dm9VgZkJ+G9Izxe0gMo882wO/7uQvXR9QFUtSnPBzoBvsBHhu+qd260b3P+k7wmQgz8XUH16hFQM
PQ7QHsYebR0uXsXEqIILzDYDsTE3YM2OKlstxZRrrhsB+0xwuaEwSWKru1l/vrislQgSmLmGiH03
udFTryzXEUPE8iYAu/Z5Q8Qyvy/8SVD6pxTWmZWX1WnD/Yd1TMTtjsJ4VtYpQlEJi6xhLHeY87rC
bSzREofhzFXzWwHLarSn64EavslEA/SWG0hrwmxBqismVD8DTueVGnD0RKeYC7M22azaYYWuKWpi
DjEEQugBH3WNYEI5TKVDe5vknXblKP79CJhTz6Gqm5KGi5w100FYup2yhYg2rG+IC5bk086Mn/pv
kPUDpcf4bI86OH4wobLNtaInK0fm/oTNwDws9DPUhYksDNGAR4R4mI1XkbzRUiuwim8tazJsB/Ji
SW9B/H4De3n9uLMidqMNeyT8fSK0Foy3GqHVCsoJhismY7fh1Rn2uAjpMXvhq/vIUR6WiC5rIYur
WBTlIZTuVddiA5/LiCoa1caIlnqLR/d4GdkUQI/W5/CFRYR9qjyhjl/uLSbgWCp7+jBpXuJCkoBL
8dgZr0RpaitGos4UbfjlpnHerRmFQ+m4vm2p6xWhBZCKTpJZggiTBZYW5X786W0GFy01wmlUrNUb
/xspoBEtCFZIb1emcKJR7W3Gn8Qd6lS6br00GsRvaK21ddHEqIs42lRauPqqJxiJDufwuTTq3eYn
Y53JdC7HWA68+Ac4gny8lNMbOC0UTMiOvW2yOJfpQmZIXwETXlD0DIkswBN1hJEgsuJ9t3DqY9UF
j8s3Nh5Sv8yai8Wnni562EtlbyT6DE/taSQEVvQaJ5swMuaFrVeipbaCPldf+erQZpci5B7QskJ3
mZmiAQpzEmsnxYbzpA/ZzD2EgirGMFc77zlN3jyCHctSnGLxRxhooIBw30HQ3sdY3mQrAPdOlFEF
e6Kcd8HxDwXDBjWVu/38P5Xp2Z72raRRWDIFZYr3A7ircoBxZOSUmeDugJYAK4OM1Sw383dfHM41
1Ke61gWs+a5fWsiqy+THMECzc2P8y+1d/zJpCrRv+pQ9n32WRKVSa+J/hCwWd+BbapXB5WjFRhIt
97HV7NXqz2VBg410r+YJZxuc6oTtKy3ADeOKjmhdYFrdORZwEZrUkeG0Une3pEzYnq5i6ey8X/7r
o06HQtcyv3bRK34Ll9ZivNfAkOii7uJjQeb353tVZCISS16hVswtCTa71RidEJ+knMZnaSjGbKS2
We+1sHoXM8vMFFshFYePj3c5j3kpVeCBFRrZmsDYP46BkrcTy/m9HDJZMg2e7t+OSYoGmt+fOOo7
teB8tQNDY3B1hEr//plcF1lqRAd9QWE6gKHgVFd7hiajVypZ1qQKoGqxGVpV4NOPhognm1vV3twE
bAEGEWWG90eOuAHNfFPun+y8PU1oaT+wY3ljCZYVuS/0rjbvnZ42eKgcq39jyDY4ZeCytMLg/jNX
80eXsx2oGltnfVFRvOEaPGhaaqkPwjdSN/L2hZmL9cRl4idwmLLoHyUukxV152QeUCXNy1qW1gIf
4CqUoxnbDrG3VP6HsCIuD+gYJskdgRSwRGLD8jVJuACk8Y6coqclmm2le/EVtRCbgJcOI6SslhFJ
gzVxKjDBwTabESbUbhkodqm/3dBsBgnCG1o4Pr5b5yE1o0i0pmv5LP96DfntFm3PtCMuSoX0n7IP
ee5D61bQg3Q27l12U+d98+p/mixePGM7BLE2DxfDD6hk0VGMPo16U6rBhDCWddW2gpO8vsYFsmCq
95Yi3qfj3j1VPKx1vAL/umgeKtJ/d1ATJdw16LESCVL0XQX/Ko/6uMhhxKTSCtqIBpqcytdTpktC
PSg05BLYnOom6znaxfKbAarjJLNokjoTetsWbNwHrurqcwoyRD8HI/j0YQvhOnGpG8Q12NVH6BAk
MDnEm7SNRl3RMzFM5IDyJFty8Itddse2XusHL8L6eS7nVCwF3MNNracucEfjMJMo1cjbaOIOfUKc
4yKAr6dj6YBdgVPmIgJDad2gkq5Bsgm+i3hdrJjGS68chT/sTjukZIlGF17Y0kCnW4T8kP4XqYFy
lQQQdOn/qasQI+pDj6Zdf7kP/G/9ijvApQobqL4rY0xdP0iVPiLsFvykpyNMGurlGUEonG6lvR2o
GG39FMOWRs8J+HJJ2pDv8Z6utZsO0D8UeRwgpE1WOwO3PYalpSC7VHaKAlC7Y/SO2qJvOY+ihXrP
mGsIVnspgw/yqLGwnHkTc4hdKpTVFz+aFhKWB84hBkeoH7Dkrdg993PV/lBmlkYVlSiXCTdW6hpB
siloY4iNKYvEzz7D6ifxklUp78P7blKmxCD12LqLFeWsfP7U7O5lDuwLRFvbbrISULizJrzKqSJT
bxa6OvPxmygzeQlTEPhYcPoYxxV8jauurIIqngpUVIF5FQ86XaHBy9Ayp1hmU4ax4iQQ7X/zl4W0
mukXaM/Hk07d1LWdtqQ843x/tEwbjGuMFDWNv0AOQqdCMgzmn921W9Cqc8lVay8T+DLvjn8E+aHd
Drnrj8D5vRsB4T4159rWoFqFLivGL2/yNPfzYCpzG/K+4fMk2nSZNn7xQJeTuEdmJSwv6suDiX5n
PQZU1LptoH3IXVkUoeHU3hKY+QVtNxyaeCgXHr5UKsRlRQKO3e0yCkf5IgiAIAxSbrdUsOCMKQYn
2Ph5TM7+aelWfA8woyMLcA+9YS5WwgUf8O6Ks6R90RJsZ4kVvNP6hCHHF75LeMfQ+Y8gtpCAuueQ
KRkSUM2CokKhC1NOARL4lkg0eSg7BnbHXDJNG/LHsSpDQ9O4RzbQFI8WmQjLq0QvUDkOElpdu5QK
2GCf6XY6xtuCp9yNTuTFUS3vZ+Jxe8qUKmNCYc+gcpnaKtP7rM6QH+0JFip0LRCsMRIwe0Kidjm8
E43u4v5F92aLvhWLlR4+iLPXG104R+2JxT8ctb07D8C5Sup7NyIcY6+1qPo3K9QUeRz3GJGigz7m
cO9r/jEW5PC3ek0Kdo527FUupeIi533/gZheq8qC4WNmGJYfAJSrKC8Foae4HbMc3CIEH/u4II1E
7TpbZKYdQBNVj5YYLkMfnbWB3y5sOE7Lqf4YOCu/7E3klcVH/LtS73dKZc4u7DiayIdopQ2VZ0+7
RjGqwmAn8YZMW6/53nKnBZQ72/FJweWTnrEQ7+Trk/+EgWPPOWFv9BgHJIzUDiSnmMmEXd54T06T
sXNr8aPZmvg8OFh09i1F9pE/SUi560PWeGJHf1mButojeAgF/G8imuavpL45/rVg7N9SyybEbTUX
YNjwXohmRErp1IntIuMzEkmeJngAsxxleB13YgJxTxT0ZlnyNdOYZjwOURr5eEpYuTptg06PyTfw
vxcm5eYLY2OvNNz2cfpCfUukunf09fEL3vEgxHfo1R3q4t6QaP2XNn/y25GQoQPWL9rKr83i5LhZ
4pxvQpIShNN/HsQ0R7LhK4VCcjYweaZ9VrvOjoCID4TDPcGvOCBQlAjfT/HK5vv4aZHM8OzwnerT
+i1lKvfDnMajD9G3C8NrRHPW+0q1JLEOVHaenkTQrwyGva7SlKR4opnlnBfi4OPz1NSO7atBUcxq
ri1KkWEK0DGMO5N023YnQCtlwO6puI4KaOckPVIiNMjNYGrQXbw5DhcH4onfwGoyvvYRdjAgRc2D
No+0uOM2LSkSxfIQRijJFYHKn4uLIP1jsETemFdNLdYCDRg1zyJTII9M4jYdYJzyIjHnGe9Xwh5P
nTPlZlQGOcrhgg05txh25v+xcdFDVaxOOufaXwa+tC2DU5CTWzzHCorUY4eqKGxFj+QUTEfq0BPA
m1W8Tm+h7ajWEDjei0lNcKhQFISrt2igNHHHyxAh0qiiQqMFGPeF9wlkkTA/hcjvvkfTVwnHsktt
IAozYqHPiIuU9zXFSFfXUDDQ+YCyssCkDNmFiLCkjfUBTLcD9a6nu3dgQuX/MHw502nmxzFIO7tK
j3+0enhF15m9oztoS+iYbC85sMQUs2WcXlp8QUXUUQVje459jpqEpyb8CRjr0T6JKmTsbbwygqYD
I5xa/90BbVWpSp1MDzATOuCEk8jSJmaDsd+cvDxWNuED9aT8a/nAkW/Tz4XnCVlOPsv7UiyB1HSQ
Y+qnK0/XrWHFwE05FRHDCZVDqLeM7Vmi5kUaw24AncrBct/frXs+HAJdhsQzdp1FJMMO8TAGhscg
1YzuE0oQw+ovnIe/gGKsGAy4Xr4XGsExqRjwqRJhlt0UrhH0ofiOOd5XFE4+gLZ0Xy+BZkbiRYeR
azZCfXsyZFiBoacx0IaChLYqeQdrG3jXh4idlUotAvvKP1i1hBooZS64B+nSwjCS4FnyjH3/Mctj
ZMSTHsIW4ofsJYJ0ThvO7mRMw/lJ44bmpzfx4cfelANfTRHr8exX0EUUsFNoVOPOWYZOom+2znnV
jQZkbSbR7WwgnYchUMKkfKkgYNCoRtwRSIs0Q9Mr0Y1y5/q7pJpjYe6XKaFf3NYPtZa8V69AuVGH
cw8UKRJW/brWO7No78jHsYpxZ/MywF76KbzIOBreNVKQ860nYS+HNo3dXaLraEmKivXTW8JA5FRe
WqEbTJvWveL/am8ecjw0zbgitxxLMKXJbNgmDuyZvQz8kXP//Obqaw16Jfuu0ktkCg4oGwuMIzD3
nRtXQ9FCsmZNfofHzOFFbCZRtqwQfU169gGBJOir9Q9bUniu4iUlK1YavV9jeL5fCyXbRWGJOqLR
QgKPzAzfLukgxhbb3+uQHhxFiBId5i1lVKhd81lGOpzmNI1y8GT4OX6Iu/TcmCVCw3AbQJRguZO1
BRG4u1hEwKlHCnal+tw+sZEHxKvu7P2YnFgF/7GFoKH+GpMuYmqGs4xCjYeb11lFpFhQGD6klMln
UchXjpkVN/K8OlVIpbBulra53ke+kBYfeDVKr5TVTjC+QYMpb501/NJq7vYC6LtjqV2JDCx9MyXu
xOQLElfWQBLZ/Yhr5Wq1mK2LrgOWDOAWXDmuiVu/zBgW1Q4zeebuGxFfFY/sQaqYqdBSB8yNLmcQ
H/dvUOeQLyTpM5Xv899sIbKfVbeE/XMgBm+uk4OgZWCyDcZjRTRcm8NUVpF6puH/ugn4LZYcQFWe
k1bLZaVXcE57gNYK4ou6y8IfQt/r6hypmT22SyB4AHTuXePxR8egKsQRGZgOXSboKlPKWC+ADhpc
fW49kWNs4fjC43tx2KjT0ge1jS46n3dEOLrep+FhzyzA84upgwI+uW9kSNSdaqOZQ6tIHH6lH4Ef
eAACUPi42dmWteUMxG/QaTOyCsWbFFtW4I9bcnxMa6NQIpvy2zBbjC96rhND0V2xqBcJmZFTH5Cl
BjZFkXktFgeM9Q1nLlYZKsYNdwMyMmUJ6I8XAOxPwwLyO45kahcbKIbKeyYU1/G2UB6yJsG24t2c
c7U7KJOxRcYrUbXQqTnqniTVDNv4izBf/MV4E5bKt8QbdAkATOCnVCUIQK85Dg4k5DPZTbbQlUK2
ppGKvOmK3bPprqa8Fx8b2v+Juo0XUps3vYJUsINsP+DgmLslcw3nR+8FZkh1VR36T+k8GqvZ1nXx
OKnxNSN5StHaLKxgncbnAlFq5di/cXzP1fxMzQZ7XYQ15fkV0iOZeT9qqGzt7a3mLUCUBRqgH8X0
j98UXJX0/FBi3pec7sCXuGk0iVeOr7JarsLe3brm5fhtSCF8Ky6dxkS2XwNjAE5GzMcA2/YWKdM1
ynJmBlFDTZ9DkkEB2vyGs5fTw47mN23WY8Y76S0VKfQlQ/YE8+SlL0U9sF/y3Hil6ETaTi8ffifr
iH9IgKp8Df4fauq+I11req/Spf4oCx4OM6g18L/n4qnhToZm23U6wCrDai8IcJ7T0vTkhCmx1hNK
orfqaUHnaxJ/Dq6bnYFrYiHQQWa7dcf18L+L+b8De5Mso12GvZENJ+emEViafxGqFjmwiUO4tnEF
aDyBfiTxSkGg0044m6/3TWEI2s1O6aKCYVPopggMfuwinisz9GFgnSIZTbrPYbj1hzClAwYH+VwM
Tc4nKbuZhD4MbbH68FJRJJbHL38FxJ/PACuhNwrrGcUKYZjtazpjtaBuJF6MAPLiiAWffUJqvUCA
sjNlGocR4RuwE6cDNRmaZS7lwXftXrTnUf+oycE8aphc9ax3brUN5lVF/AfIzlbBP2ZwzsQ0kzUc
yESIdfbP0Q/pdAwz6UvgCgDGmaT9EKKfNVpixdsc5GE3d10AQcehgMrLytFB/J4p5wmWm27K+ozO
TaJImS04H8mu/gWoaFQUoyhVfJeJIiWB8PWlTsnlBU0HQOJF2wxvnyuTaGIQJODgf69vbRIkFM9H
lXUR5KQUtZW5wh44QUsJbWhuR3OXNRlnO9A2hw4GAr1JjnYWSV5HAs/8xVtfOwJC7Y4K+LDQX+Mn
z+DaoO6hxy+a0U9DHd8vQX1G3eQhN9Fz+QudoQbnkGh+2DP02hIvCSWK8snMVlP+n1YITsg5zi/W
WGWaFLn+lDjM01O3dLNvV6TvYC6O4fMxyQKpQ0AmzEAqcXsz54PSJcwA4NJb9b+6MDYwmsnEsJJg
s/L9NJQUYgZDWkyQtMj82Dd9JCiKfO38fYn/YcR7kU5JAuHdaPdZACnL4nLkZp9KrWLKcJUWdUUQ
pUaw58BxqlLteBggloyofobNrtLBnbj+0RAimlTapzvmOYR1qMqJFHSakFXAr5xIRzXCwvNKuO+S
r53u0195l+cxme5AZWSJVYM31Py+6llGorr/swT2sOUHrl06brr0aUvimSs6PXp/j/EtvpQhlvkO
I7NfYcOhoTQ4g+0moTE4X3y0NpQ6mfFyAvKk7HTDDl5pcCPUEZf5zwUXckf0oHXrjzXAP+kmevME
65peYSGQckpPhhzAsZC2AmJ+lWkABDCDl1t4rk89DwO91N6g7ZA5bulOJOBcVQ7Tj1XWQqnonjKd
v3Awc2UAcvAZLcNuJmIu8PtkL0Wp0SKoPYnXHDVZJt7cJ/eHUcTgWf/7MMbHJjFM1/W7larn6ym4
27Y56s/VTPgtq+Jq7FHnMuasKVQPIRcfGkAc8BuspEQAY2jC8cmiI9AO/4BkHaQygOzqjPIHOqNz
ONvBhiLPP0sXfkE/ZUo4qM9Vyju3ayIOzgdLgHmJGUH1MVdSM43VY/EVshppZGh/4zsNVw4LmAay
UQy6r+arBoEtG5jSos+vJ6102xgQ7Z9hhk8dvWiP4W7JQNgRL5wInip62vAPRr14+FVO6CE1kJbW
PsLm3oZFi6Fzocm1eEycs48tdM4K3uCx9inNAYZRgWh2mwz5/u60Lr0OKSTymceHJl/sI1UU84AB
/SqJqB/ektnBcA7x2Lh0XeblO1XhwC7ufmlm3RMDlm2x798V0fzfrzD6vkApLJfoW0B0T7JELS/l
zY3Y6my7lh9hK0xc5UIsa8lz+R9Dt4IEyU956CgyjbhWedP6gAdXxxI24ckvjkmnn3sfYNQnkryP
FsYnrzVtIUSqu36bO8vlRKtA+sHRFyhzVmJcVD1js5VERIB83RSMo51I+gFyuFT6vMqmjWXnyb1b
NVEo90pWHAFOP8dc9Q+7IrTKuBorSuG1kfGhVXemPV92e6R/IfJhn8P3KpfWuClK0cdZMp9Dxfq2
myCpsFnQ9T0twiPsrvM1IlwPlmtmAHkcq1FpJmeyroqbo9ZZ7ig7hNhRAkMibKP4CQHsXOCUMR8X
ULllqmGr2IPYSOqFzsTFcFi7yVNxcsAf/ZddM8u4FuHRX1R8zIhII25R6l5CxQIRTuGYz72YGLid
SHt6Rb5jCuAVDNAMf+NSd+3JUkOOUBuYPc8WORUl3kSQXi420yeywX+RqZyN+K5nhQjDHnsGqE5r
hM2QSohN4CQEeAeNSAw7usd96Eb0pU2lsZ3s60sydq1RkjsjK1EfnpD4hdF0zotm6xn9qcD7zQTd
0GrwRcJX/zbIYR5zF8lqlC102+vYr61d6VA0u87sUbZD6O2+3SSNdS014ca5RpvhuU4xMAIKdxGd
PWDPH89G6tl60kYOszYB/Im3USVHTG7UpJ69SBKZd59j4VgnMNzL4iYbRQaZYmrDKbu9NIG4MMFM
k1UqwDpuMI2DSGoA5N7+NNEdunZf5ceRZPUGShls87CKmr3NTHpYUKjb1unSCMtRe08Ny8zSDCfA
SwbafI3npeln/Mjbq41UUKkRcQW4lh8NxqwPXM8Ez+h8H7w6XCw6+dCiWSdqqJxFojr3R6sChYyB
NrRByJv1D/3Ofqw2lf/ObY5khvasVBoMGrjyFb2lU1+WjZuJ9gXzUgu1GkG0rFwJYYvpT1Y3Ux1Q
IDUV5DUFD6HtosF4+QWdVF+TUzLEEbaXenDzizHMjPu3GOmiPmkkKz4EUPnvOccTBy9bFpebukcD
72TWreap+Dq1xeiqL1PLcW6kY4HCL2/ZjcMisOG2KCQiQAIXEp81xioc97tA63ICX0jf0/chyIMY
jrhPIEIOoR325Bp4EHCJKboYUBEJvZ4RE/YOJik0VB1bTdAoZQoYpoOOU98a6cruQfNNR30MZhmr
Ee7bt3yJXlYUET9LHD/4DHEXkgcc2Vj7v0NtdP9tUfXSPYYz2mWYV80wXlA/K0ZtMSw6IZcj1+xv
4W3s+z3eYGYJx+K0nBhpYAcpNFWs2R5UXKCE3xgEWTzZyUiBJFooFlcplxz1DBgK6hZApd7WejXW
r5D6Iih7Tfe+aLLLqQj7qcBm8uT2fF+kFb87FW46W0P/+qwKuRjZF/2PVCf3BA6F3S25naNvrGvR
j9eeUoPFzZ1X0hMiq93doaWjBl5RelexYvn8azJ3ZX09E01MGg3QPvKP0A9f3A6r4bq7G8C5Eykz
x5pdjqKWWwVyA84mMz32/JSv5B8H8e6fAK+jA7tll0L/jHXArO3clzB7bX12JevNlEe4aoj1NjR9
UG/F76D82g3W8VHKm9V/JQsYqV1TVY1h/g8cAPCAQ7z89ocPCz39+t5nPvqPsaV98gkddPQy7cDt
VRDu6OtczpX/fCTfNRZsaTi+52LGp/UpFH20HfxVj9Z0+q/9YzG5Kk/lgm6RqC3P6pv/+ubRsXNX
p02X+V2JrSVrvNqkEdMGMKAQ8k0bJuz44TnyS+kSos0yrxqdvNTKrtb/CdxsEpCnOjVVxSkolPhD
S32F1g1DnpibSmGrIdX4w40TEQa4MrfriUrCKG1TJDl0nEqYE0m5P+RCjCQSz+Yi7JCboX6wewwC
+S14n6EZDwHk9Mju8oiFeSQhPdxl6s2m6REby60BDVwMiUgOe2UDXYDduoNUxieJBsI4G8CIlI8N
qXCOt+Kh0Z6zOAyX4cOVgamn9we7Tq/0V40C1kRI9cXz3t3wlWcahoKSkBkONNXDJLOHQYRWiU/X
jwM0DYBCT+V1M04HDWakEwCzEFklGwaHvUSswbdBJmkHduIJRY+1fhnD54nDGsXwTNXotppf1403
zl/i2cDlzdoXjcq0xjlZ3z031CE9njBTVrDuc+OrEiQZGwSPmtQ6v4h7G+6DaNdl00uQUGycG/MS
yRaO3Mh/vqdGE3YgcfZxoUnuZYzTL0ELIO6CFQo5C0giaWZ6GI22sSJxMzcLaJJ/HkQPe66FEklD
+B3zjAIaSGlCkjOJuH+fVa1DTyxZo5/F7mBaHrmw8k4XWRyjhqhlLZ7zbS6K+eBzCm82omwuNFg6
RDbKpLo9PLjXD2Xju5PtpWiiRANcyeeHCN9mQirFySMtGDW1QH3NnPeZTs+Ca2+Vd4YxdCysYRAU
KDjr8Qy5sx/V7FvwXrHgLmXscYIU4ujlbVNHEzuSDZ0MUwb1aXL1mmQI87Dx2id2R1Y8N8tUc8fP
8OzM0sx3juYdpAxpQuKYODkxvEzFW2DG9QoMXAzPHlBEEC1SinFBTGPGBDB8yFdN3/LpE+nou2GD
mFDIUaLNZLXMjRQdPPs5NxX4ggwC0pBuOcjEYIq/Kb0q/T2+SQXtKycRZxZONuEiulESTNIhCoi6
ZkXXXumUwafMgD1Fbs2zwHID7iVJUGVzZG7JReN/9vcdTRvzjf0k0CfRZc9I447EVBPTvYTUoY5G
HWTLuC68cpD/R2YifBsSfYngrD4YhG+b3inwR8KUA2QicykKa4HRDuCPUvzbZHDh3hzfZk+zcCBf
VstO3gp/xIoAmPT1H6TZzzfzxEkA1ZcXmEzOvl7D2FrHnJRce2HhJHw+Ah+9J6teJgF7LRJXZUZe
6iX7kKcQbCX5bXHJpK6uBFnbs24bdKcOh/8IdQwlebXysJxhTOtSzK78yedTrc/otQ4XwWZ+hiNN
Fx0jPhMKzYU6fyLYewfKmN1v7izBKNUA6RW2dJGtMQVTr5Dn4ueoATpqJbeBoxLGVIQjqTGY/G7Z
Iq98dOf+Lh5vZr5w6BPfFEIP8sXfFrMDpro5mO7On2NSy8BZMKDpAKtwqx9jt4X2jhcLbxL8FVbR
a58ui1vx8OWV68ihomkSL7ZjMtxeKIqCmF9NR2aS1JA3Z1SOtgdSVfhCNat8OdaocnD4USO9ESJ1
lTNk+CbiCg2aeEHV4L66hn/O09HaIlF5oiXaTIonqdn87nTYEvDz31opUVBn6IIIxQYB2n0H9+AB
rAbrQodt+6NIfpnRJFrWNCgY4ngBpH3JrmcCu+638QMqJsqqmXHrtONMaKJRY2CSbqLj5PGjSRkg
BclBlOnVLhSA2NKT2nM4AfIJ1TXJPURWHOqvWILA9K6Xhl83qfZmxzBfPaPD5lQ+cRdwYdXjKY+G
wVsGKJPzxgm+Cz4CZuWn6rt/aXP/Y6UN4/XPJ+k+ULVj/+lGLT0mpNO4ZL0+qhbqIVExpQvI3nFG
UevE2RHHGlDEMOFbKxYJ4A8cj2x4TW5+hRYbmZr6qxl3+OCB2FcDmx1W+lbB6cZh+PrIamRtqmjf
9yVIPjRX3eMmLJXvvuVpwzxxgdYIW045AYHWYg7ra9tBsaoen6aD4C5s7lccsD/67IGZyttICail
//XRQNzJIA6WecrMPWj9ycbAp3Mg34BgylSyE4FP/dKhTFLVmYnKH/uwYvU42qVedejNr6KtLePC
bVXuF8Q1ZLbSfBuBh0Kq3Zb+F03OPCR5hkHil6b08IZpz4moFQfOFhPnq5PKuJ7d9qZGwRby2riq
VJ7UBRPHI7WfupaTRkDP3xsHMpCgDFx0csKCEp++Qti5T9mHHHanAsaY6Dt8tHvd8bC4PQ5Ay8Sg
/M+pwnmmAUh0rMIiegVFwsxzZcy3bdLDZFcqFGJo8cIjQEglTAQcp+qLtcWlgfy6jO/0/bWuZ/iE
6TB+wHFGEWomW6XZpnL6FfBjC6SI3tQWjVABiLIs7LTjEgZVpKuShAQZ9Cn4e/Ijjlc+bOXdZek/
Q3iGcvGsKQgUVORtfx8S7ASlqBJnNG6NYhRwPXmrIv+8bIDdj6gP5hqkLMCY+9UJt5KCygjqPEKg
VSSfZ4HoKkmGuYt67F2vEEhSaU9qeQcfavNaRc1D1HNLOukqtnzhnT2wQ4TO5AcoviXAfmlJsoM6
8dTZIUSoris8YghxCxolXgmkuNov9bUq+nTpMg3p7Sz2sOxWSfS3X93gt0bUMEMBF6OwAZwxqmef
c7O3FnuJFimvunO2qtDEMBRJlXq2B1Jv4AWz88QZZqoLzR8WWoFm8/u/x0erEQN4s42x/kBL0HGc
bdIIYTYj+SQXzEsn5LdslYAyUEmw4kRBs0uA4lu0gpMCBZxtxC1CN6pDjFEU37l6ES02kIbEgPT5
onYeiSiK1kGVLgT+Dv+v6loPEq+LjI+FtFHHUasimJjcyVj8mc6Pnpo0/DWouVhvNklsJ2Q9o7xi
NH56BkIVjoqQ93ucPV+8nt5/IoLmhsZY0p8bzmyp2oDfQWTvwy9boUMI4xs+MgNJddtuA9KbYBI1
PsWWYbsg4RGYfsldurs3NSx1S7yi4BFOmEbU7xNTxGe6zI6mrhRCZqJvaYqkaCJPU1PWMYWnF8i9
t2ct8jXFxYKVdAoDH1cK2HKnhQOJ8H0nufTZlfYeRzrkWQovm96pOGsvNf/b8j/2zpC/obT3CP2x
/p5r9FTJWbr4kuqvZ6yRo5GwsGjtsFWFIDngELTigA5iOVarJy5DtBFlfEHLyOUoycOSab53i9rh
QEf1+oo+Ma10Sr/D0POpuo6rRmxXd75NxhcvZU1h9spsiBKCrAZuwhpS1c1LFtxOG8i2ijf8WL9d
pD6SrRS7iwLunOXj4Dz2RJLAq5DpoOXQRqNIHXuGmgyydDKCcngDXryJqTdvvCkgouEYKEe9R6ih
7JGn5TC1qJ7iNIGomd1+pDB/uYdj/9ody97Hj+usFzr4yicbdweyJGwbgBgrU+Sz9gCwEOMdbjm5
622jxHeAobFhFOH3ibZtxfhBOtcObBlrq/kRFB9/3w25ek5aeRfJ5Ku4Jhze/FiKyORAWsyw/C7Y
GndzqzSu3HbJuFAWrGCYmFhkWHksEiX9Nf7IVPlnxhN9q5kDBpfa/4vEZ1IR0rk6ya0JyVLlz1OC
dL6Jiqt3Wacr8u7idNaFG8syTlq1iMWVH03lZCiNRoEtx0Hc7Vihxuj5MK+HC1luXR+wNAwqwPmJ
AP2ovGlsINuaBIOEdpXPkVnkjCiQhnNjP9E0UfkngE1XsAn8FB8vIC8UjTV8BHCJT/4HyJ3wijxF
bQrN9o6Y4u85VLYjj96dcZQuwyMDKMCiR9cbNrhKoZ9k1HZmxZJpOSJNKGC4Bs1SufToPuu7ueKv
0dobIF5oHvJ1TaGROW+4E8fyPCZaCr5JJuYIkB4tZ0fMsgQ+2zz5rKZt3bew/9Tp4Dp7/FbPBQ3e
eyn4hPxkO7HTlOQj3MGBpPLZ08++21L7gCoh6dxLZMNhZCRb/LTU+r00yR9V0rBDMF/fDxBnOEvx
MRDxOXMrC1ffS2xJxmLoLae+SFScMnS5GultY97LpEuxz7oleuB480xDJKs+DhTDDGZ57TeoOUpk
0vqLQ3gUrGYlanxrl3dWm9svpopxiYqYHw4o8lFdi/kOxzBCHFR/R/QGthRkgSwaEHNSDK3ZtVmJ
NU8rRwiR4DMNJCdhfs+171Y+18/jFjLuU4zobHY8CR6Kf1mT50g1VVL05F66+9QqPz7ZtOvc/QBc
vb95ESEE2JrhHQIySv5136LI13py79QjyZIgir+en6POjTkVB/Y6AEri4QsIyUuGqmfNy8TM3FWL
Lxot+oziiRAw03gdXnfGde7HO0XzV5N4OUxQ6gzhSVoFYthQ0kqa+WvdpymjTt2KoY2+f8sf9bIq
0+9mfqT7xbRy8+CcTdIhuMiS4jGu+gCOqtRmFT7CFuE1OHG2AQn8HsvuBO0rKNnV9JBo14cm6+hK
Ntl8Tf83GqBbFMGGS0KCHRY1AnTh522+b6vuEj9XkvqXv8gSSe+InvzTEtKFwz6rDo+AdAajWI1+
3KThd/t/pmu3IE3+JRMHoCea+auThtVEuwkvi+Y0Ic1azwj4U++C1E+4VxI4DjcnuX2w85GhcapX
diUU7G+ih7v0Ysb382GHMQU2duIM2axfbuQ4yQLvSMv1CnoHLSRuErR11+sK1nGgUxVEUq2Qv4Wq
pm1p2LAMUIP8vCUQ746fFMjLioRIDaGT0UhwH6qV+elQTbWn6HWTNgYL4n1zI/hG0jpxbBGuVSFD
KrzADE3K61b1wuiKTqFpPT3MYsDaYCqolbSKdi7RlYfPCykV6gbfoFDlVYoLimvK5XyEI7h29+/x
QqetzZ/d03XZkQ35M6KX8BZIX1SqZnAPrCP7Z2vuo2RzTzu3wPvWNLXxHMUkTf5vs71a0+Yvg5ws
tk+3BsiY5NXC4jfTyRVtHD54lFmrxLYl8WzPZqT0jmrFAnIwb2mmJ1owPlQHPYFvc7gTzygXEan8
z8a9mcwxZ1wNy9w1LrjRsR2eSYIGpCh/Mfbu0HKKjj3OU7h5tW/c8FoTplYsc2Z7d7FNFuYdrCI/
4GT9Yv30xW+FFRePZp3R6DtAktsORTKkMeIEGyy7xbblcHtuAXJElaAeSbOeye/6+b1J94qbiaSB
ACdK+jgO2SQ+IyRBwpxBx6eTf0NJNX5S/eGBfPtrx/gIRxCDZ+NBw9hI9UP3bjk8o81lLE9r6zpu
sgNg8RBqiuxmI9nrT87++zrR6WvcBf/Zz+k+GwEacQz0CfyIyH0K3Fu/yaUt1J4Tzzx6SR0mXK+i
Qa9JHKUR+9w3v/ajUhNYrfavN3A53HPEwl/yo7twRVdnKLsM1TBgA7HH1czChV8GdVb5E9oxnIr1
KPo15xgyLcmQ2+IN4OWsq+nCX8bNa1plMPLcjWS0HYMnS7Fs4pO8k8UFL+XGnxadLuLJoz41p2NA
tAmdZlCV32OVm//Yh3bm/kUEUtO54VPX1oNc71sjwXNnUIAMn8tnYwthB0jYSOhc89Q9B7CgXeEH
i8aNcDWXd0W551o7YwlCU84mxB2NRCk2cDJitibRuJc1Mgi9ttgV/1/1xofZiXyNwVPJ3Wf0UO60
3y7PaaVAlUiD7QJMALw2r0CjEdrPLKvFxAHvZ8mrAn/EigGEBaLvkPie+NDKkjOePULoBWA0cclC
06PQV6kL/Op1j7ZQYC0oSAmA5WQDHjyhT2fzg06Mt+pgRxUEx/lGRUAc+hA9iwB05/va4Um8yPsQ
w7yic+1tFT/ssrv5JSoZ4mAsP64qw/VlmaHHNl7VX5T58y2L5H7a7yQ69Fladj4/ipbPPkH3rNHH
9ds4DTKkQFudWnl+LHj2WepczHsgsutXJ/KnmlpQszmpFJdBvGWLQ5yJfjvk+EOC1Egs1SlZeOpK
QM9To5WX9fuoOf+6TZhRYvqwJ2MG4z9DN34gzLfAfJ9eUtza62IV/3rvEoZfoc87EXsBIffMqizw
4GyLRqjmLhsyUmK0SB1NfN/UlvW2xY03L4v9D/sisyMFWMlOWN0xdfLTAh+yoZseJG1BSRL46A+A
uSut7X+TgoDlvtVCWSMLhDlenAdKlN+xAd/TtByNnJgCfaaIYSjSjWAf2Bnw8JxdhKyMNrgo6ffZ
C2aTRli4r+ZZVZCD5IhX/1oG7/RxyXodCC1oyz9mNbLfVpfJq8CzauSWRz20vsqvbTq3VBB7NmQC
aAWlcPqd14n6IqY9ieTRWojbiCTjDnyu6StKte7AtpjYR1wNws3vXbkeV6AHuAaIvkm57cHEWI4I
9j0sSVHk4YKWZt2akSQBw/a+E83rFlkyxx8ax5ixKftDJHbFUqAwcPyTwSG/+wIxsVEdeQKsuj0F
IYVKmpuTbLN4dL5lwcTa1qg04IdDEU7NB9lOyjDZPLvBdkAK29rLFnHIu5uW6rXkM4vdMquq65vc
ayLcnm7o0u6mIl6Htqx4vNNEdsLHPEqaOfL0N341MYzddlubXcFUC4whWxYJcHME8lcr4rYudJZL
JmnJXsKSLbBQLIST48eydHG7tOZJuFrNUeDsnNXSvqOhMt4PKLFD9f5yV3FGDsLLuP7G56YXb/44
s87cI4lDPHJLaCUm/0+F8a++CdOCX5nkg2qdtqxyo+fc690jYr3i5d/XVDY0VpJqWx4MPB0kIluI
lDUL7gUtJ38vrzfjigDjqBNM4k2VUyHDwkyWSnOYSTVbQEfAZNI9Ocf+E3wWjYnNz9qXby0FhvIg
YL3Y0R6pVG1ZP4KtheVxtNhyl10tuLNq6pkj0f7KMrptxRSsH0X6yMZB2UTIK+/Aq1FDGiVkZt94
jF525kwbJ0C8qmXZ9LubIsBm3D69czB8T3bwBoXFFuA0PtVr6nC0xxMVtgEbg4YgDf50jkS2oUVO
G4uwIDuVWixio+XY9AqwL9PlNEaH/pshx4jJ/ggcHgYnX4rfkhudz+xLjyrOtL0tKG2bs80Zzw5+
0VDSX400bitJ7ir3u1UMk6T6vVcLCZo+Y1UAvyAhOsudB32h89FQCnbQ5Xn84ASLG2AlLxgc1UmG
/eB81eJe7I6HMaVhEdTu22zaI7T6pJsVcw6YFB0km1kZEualOo/rNA2yVzavpjlGAAzJ3ifAX1Zh
Qwvns5rJD4JJid15MXkEBewGVBJt1KbyxbGTpR/6yJPCzO/rKKe87xGYVfFjjVl9B+/ysRnkJkZ1
ryaaTm/QibKbKeBR3IMuFBhLFPjd0em8Kb81V1xIu+unbLJeu/6Py/nVegXzknJv2Z3x6kBzjDSI
p8EQrGJAP/SQyZ660WalItBoscoog/ISXM8SH5acPXTJUPeCJ3LZUon8A10ywocFWj6GV5gc/xAN
z2VRbqYL3lbDUJoOBvXyQazKl1DIAgAkOiXBzKlX34UNb3GOB4f1UOLc7wKP1qiaqqzPy51H+AW/
lRNisNtjxrAV2PbYL8MJXqK9PNRKHuH7NAxL123oGuwxDrrhy8FoIa2fmH0F23Rn51Tot2spdA4e
Ncfm+N5yySgTjxyMS5ZnBufTnhwYMidsm5bhPX5yjbjLL9IRunlCrqWLgtMGihxIbj7VfUOInNz4
aGF681EjRkjNejV13V0t5TdgKkaK0QnrTFxAoxJNKW03n3h+J7g84vtfsayY8heOps/1vzFicqfG
WSMBSnf4skX69KNa23y5fBqMy/Iq9KpKzbvRpLUKA2Z0vAv3Lv+LmZQiGmaI/YOgKkSKHvFJD0Hl
AYg5vISW6HpkLVE5slDb6IG97Ml7r5w+hdg0QYvWbGzbee1tE6ukXqgD8nif/3qDekAqvSe7l3YM
h3GFy+4xugmC9eOfpTpGdXsT0E/fvUsMZRrct4rf9BMh9qH+/RxqY8Bn5bOvTkGnEjpowz7rGaZs
7YahA7a+rzcCQGVT0TDZ5Ww6SQFS4PwTIQDx/8SX1+T6PB1oauVEbfPrV/3Y05dfE6sSoInvIt22
kxNDhOKcLdi47s4U1EJJUN7PIniIB2E4cfnNmJugWCrpYi1Hf/HVpDaT37l49dtBuDYaxkZYgQPv
cKhf2N/6f8cvo20V62DoJC58XTQWpoYDVfWGT5Z8Fcya7kViyIm7sVLI01WQWecm3tlKmsokbtxC
mtFO6eEzZla7ZV6NbizpaFS8yPzoPnXdnGRuqfKLAzPVTzGFAUhfaBLLAsIrhvNnqu07NA37q9B2
e0bLzNPxnPw/0aKQiSlw9sK/Wh1QTlWCZIE1iDO8fpZWbwHMmsiRUSJPeHGbsHXOg0kk6+HnTAT5
txH61feSAY59Pgofa5bY2eq/hfBRXOwb3IWY1V6EvJsjpBZYLYiDf1NDXy1oteFP6XxyrckUQx5e
+Df66zKIt+i1zmld0iMrHFq84c7NLHiP79Jvx22yDJwlGiHVjnP5/m5I7R1Sw4CHOf5eHvqa2VBl
3w12aL9GtQsXGShlM2FiYfrJhQ3Ldr6RpHKk9MdRoDs+vbdfv3ojXnja6PfiqpxfNm2FFPvRUJHB
mTrkOwIp+7Ga/51erhW0on8z0MDCj6MbEtCNbkkDE9lkDuZrYUXUnirn/iOWl4mgX6tEZnhtbFQB
hjixCz1qJKRZI/tlOQyvirHn76XMpd0VfNbYCdLDjgao/ytjRL/bZKOZT0FNp+F7StrxUJ2MPGjM
0nmrH8mC+71I6WOU/rk+iPUbHXr0JkAVeWq56kJvLQZs8JcfF1nicq8aMD0/+8mN0HvV7uY7VJwQ
ENrhXup1kAb3sDNcl0meFIbGxRmK2Vd7jqLFDJcbFlpqBTOGvDvBihMpWJwZiiwssqODXBmyIQgu
mgzv8aBswQb4B9FrvywcKqfPmd8tIyzwi5dj3UW2cramOwKPRyJK6RACVWJVnjNdcx1SlsKZ3b2g
yDZtHzfXZrLXGvRubX+t9y3cuohNukssi7mTUcH9wPAUi/m8mjU85cxatXTbLAnFa++D2V6bnzSI
FvU+4S5sLv9vKEQAKcmSRNOb48ntwvf4qgrXO8hC7kwOOh6sICxmupxzmL2Bph46IhJY1P7V92go
ynvjAKEBDx9sRp14lTR0a8X3g5eeqE7R266/Inof8yT5z8el2SDE9TNI1w15dX99nVAUedPOUmnI
p8f/FkrLyYhYkRoCXEpmaYkSCjsTEQGKg6hjRipBBZ0IqjOXzCF+NRTyx+CzGZW8HxRiboDvbghW
ry1TKi09fUyJRYQc61R8cxT96pQSxJkFSRO6ChElOyzhn+clwmh0lkkjKIyxJr2d4D45IPBEvokd
K3ptjduybmlS009gslrNsCFwJHntAy2Xf4x2GB4qvFktJUaHywbbHEaekPp4Lfk8/+bGOlXRPx2l
balB4Ql+GhiViBmPjrQfVBeSOEnbY4NEI0SL69bPs39Z2VgGmlSfDo12Eo32nTfLr5kLJQG8vSI7
DOJZRjZ5zXJlEDLpRiYox6/lCpf6MWlYru9ADvq+FaD4Ig0Jbn/sYeYqUPhr8U4gepPHCpTJe+Bj
J9BAHA7J3TWRbA/a2b01f5dpjaM2kXjsbLooXdr6KVWoa6smiSKrmKtzNA2ADU9+ZjdR8Wj3gb/d
mJA+QcjaTI1aYko4aTpQ86DZ2O5Px7hms4/tOVNSyWfc/HRgsDNIBZt4RqMVI4J1E2ty4bBtDQWp
ysmGjo1L8CxKsxlkYc/06lDoWIMz/plKM5M6qzVDCKJFSuGSU69Ee0AnVHztZrpqDPk/w35wkc42
ZehdUX2lhIGg3c9PGsolafFsJD6hHxkKdIJAA09wQ1MI3QvkQS21RV5KxDEBXwKaW1s2r69Ska4C
yUkOlzV6h37AHjfM+jBp1JDiwLtxx6br4kysX6Pv29cKaVWgktPuHIbZ7qezU+pvmV8xJoi8Llb1
NH5Uu0r+Vul50RxZ81+J9jCt3N3OGm8MQ6jF3pnFhU2AYtVLcBkTKLYYR5fyjXq2kIupiAF+CGzN
EwYZ8i/QmvVXxVCIcveUMTptvKULpvZQhxj5g0iyhL3HiiytXls+yeyLaKn1bMdqQZi7+9fWmSYR
V06yv8S+a/1iyEgofrz73ifrfZO+EAzHaE9XzCkEhE/6JPkjXZoMW/4Zx6/o58l7EP1/ywVKAB6K
7cie7h64mjSmMJX67DiCviKjCrIzTrf3cjz3j+NTIjsrdg/xj9VSmIe0sPb1YOfTQ8NhL2PE8jse
ZEk0ZM2lVTznCLcN83xhCUFAVj4jTlJdB7PrjCT4qn1QxeV6cdZc00VO0OZFv+3fi+tld5ITaz6X
zkWu+ShaZQttI70U7S5vBQ6Md7ePBbCAKV7teqx9tCPfzQekImNXmN+sjOGKlZSUnrns0hGROGEf
Rgkj3OJtrXTDRWqYKflkLP66TwKfEGZ5fP9qKPS4AietEdXkT1UW95ZM+URpurZC08OMotFRvOX4
1g7q2379rZGwz8asKHM+nPd1nQnzrVbty1QNJ+Sl9hz/CfdUMHZhnv6KPkfWXsco/xq3pDhjiq0K
1wKfJ9cBeQb3+YzNIbUrQ4TLW8jtJG9751xozQHgprO3hH7xPq44Dejr6OIHQ+uwINWHSrAuRlsP
FTTCBVo0uSa4ZDyw8Cq6ZgVgD3uJ7VlM80N5ouRShaP7bGdOHyRTZ5B4ekH+mF0islz3XlFymWFo
r9PJ8e2vJ+SsRDfi5yw0zEOZB6p7Rk18U+tT11GXknU5jGh5VGswg1G0Pbbsco0kxazlLQWI+qR6
lZ8+n/MMLdebERfu6c3lmTzHpU0pAeKPmb/zYM4dm5Z9wc9oMGk7/yGT1vB0z7OJgIYy2V0wzJ9+
+b/qWUqJuH2oyGsJXvyT4c2v+FBb+5/gCT2LnmmdHfD0/wh4GL7BRJCaWgsK+Ox8qL/fOu2N6e4X
lghZJIe7e78VNJQJIxJxP8OwMQGPCXtYibDNqnZcxW4IMp0+tV2Ohgcduk3/qVR1aIMKKoSKjRYp
q8W/IWipy4cfFCo29PCw9YXRQoRVIIeoWj4FEpZPtv/YTUC7DQyxqtjGJLNkW3Y5V4UxJK0Sb27F
LpWoOsAgl33d9i0ezVwnX1x1k1go+BfYEC6fpFGlv8d9XWXtp21f3vXxUcE0agqo5EJuiuZq6oqg
UhLO52cURML2MvJlOTEDYKmll7m3MtI/9GBiCtPoXaxQ4Yrjg8zOm9Wiwd7gyblvcvZST10SxciX
UFt6W/6/sa7fX0I2Ki8DEeAW/BTxAJvut0hqME11ci6vI1tLI7xsu3jmUsCEMslDB19T5i9lZpa3
5/ZJmT4EnYglt+qGso/Yzpg27SewWGDVJMxaQFrJjT1anPeKkTil3xL0TX2gkdrW9xJMjNEssGDF
jh3H0Z4FmPPPi5+ONS0pUwVPK2TemH/Re4FQx8FN2M4ZrharJB1QoqDRJstk+7XZVVnzxXRN6nuI
uHfmGiRmfFvTrqbkinAKEK6e0dzh/7Bs13X7kY/x5R9i0hA+gfxQmc94HihTgmXxLDXwkW2/mR1J
ZSG3cdoUTr1CWIh0HBZuIb1DYDSLOw0EhSbqHMJRxp27MFRWvvwPv7kvRcuwkXdsPZ2fSENU4M6p
5OO8btshqU3EYGcxd2GcgX8+G0uhhm/KjoLpyWLv+1/mCfF7TxYJOeIYY6JIEkmqN+TqC+RNnQFo
mbvuzgWlJgHEue6bgvwFWoGFl9o+xAeEuubeschaEmdC/Rr9H5NSrk53tTff0FNClWsDr2c1vGWG
0XxToWWGfdpDti9Rn2mq+aIlnGGkunnOLQEseODtXcvOYITAYDR8fEptOA56LDM9+XP1OyMQjR77
D01ZoSFCJMg752JMZ6nNEtiXnuynqAElVV8fuWhxtaqfgbo6e1eDxhsUwNLbvhVP7g5jeTmFnoAw
/Nxh9PMrDf7yU9MbHxiDAIIhX7B64DQh7TdngOqAKHDO5L6ki8PGtTUyd168gUZuWCMIJoFhKny4
1WPspgrgfub4aEFl8a2tU0PGIregO2IS6L5SZdqSGrG2ptPwWMwxTpWyZboQRgbZWWKmpMkrcqa2
kFMSRvcwBMkEsHIirAm6KSgn3sHeQgQc5a45JcNxUgc07JvG72+emkeSkHX64L2VfaIhXId9My/a
l1mXT7RrsQQkxXVbRMDbUc6iYuX0iPDE+wgB4//buD6RoMPXiKG+TDaZ1PHmYfYmtUG1qADRPpfn
PfbLJ/Q3PNRqGmXHo8VwkX4fI/pW+rtj0Yol/l+CBaNfcfdm7fvZXq87UlN6BGQwvAXBfkvsLNP4
tJBtufrDmNf+0jq9k0eeg5Prs0sUhkkVUGnR3EtSlQOJj/G+3VrjH2ufCHwro60Ou/y3NO8YcEcZ
xtW0yyUf4XPZELlgehq1+1QRHc7QEKfypRwtP+h5vYUplIyJhQuFjLAbLmGktPtckegSIRMY9zCR
83W4dubk+oLpheRCXhn+r00jcN7AezFY507c/8toJjUjAJnTTcfgJUDlU4NKwtVPW6IOe1J29zlC
nqtXt8Wn78dRgu1Jb+s47LSQvKvZ/np1E491Pip8cbRSzIBVQupq+pqr37sTQjJ7oWyryf2pvwZt
YDIvLihVeMASoEJBwMhbGFzL33AznjI+H+0hsYaNH0Wrq+W2u/r1ItfDwo1SkmfPSnhsXkk1BUfo
RfB+FRB/53Zle4ApxsTyqNchl96d5QNQohRCfYDfWOD4aENS+wCNhOZxKG4bDwKjIEGN4wiPL+Qa
k2B+G3nugYJfU0bzDq4UtmUrFwem6lOEEy095CeaVoV/ro9N6FHtcP6J0/fjREfwIZfZZ9+F30zc
XyZho+n4y9HICMkZwVjrl6XDcRdlurVAARhUhZ2/dJUp8FXx6xfxTnn4i6sNwDOS7Z+y40fiDv8f
NqYEbNi6L4+1P0eQEAVzK8JoWiqkhG7bj/79izcgue/7OJ5ZB91nkLvb/9I5urAtiSatINWJBpXV
BOozpjAOxKzUY0mtJxLCi9wf4gM8g8Y7SGJi27iH+sH4Pi7g++2hLgevWggzroGZ9ClcMbVX5wf8
C8fGz0xXY5hHoYXSKxtz1BmdO0J7+toQQiioSXUu7r4nEJTPLl+zXD6HhnqOun5zeD/LsTTiTkWe
mGKnQeDPbSEiztqVFuGaZSYHS5mKmhPnjBabJ0WGXSdiIk5M65y2/xbPJlRFX1YbOcWv4+4bbXqy
VEsPqCDgOsXwiyKXbAiavEsGqPo4ZaSC09rA2AKHbLtipjX1u4/sIw+//y+VztIZorht50UyonSQ
BEAFZk1qNmPhUa6gFbxR2VqUuL09fLYlFwremQAmLbMedk9cxiJbk0gBhcMu1/GUOIgt42Ze08Jg
1BgflQ0//oIkCKsAMMsz7y49fUIVuchiiwUA2DplGabEkOAGJRGPPfcgCU1tnAguSsgVAdAzueEE
YX86BAAudR/RgTRio9Zj5RoYIHnAv1WiZcff8w5cTcIumOBLKn6lroQHMkfCCNuLIsKpXtoB4Ab4
W2JLJ9CMXRepaSm7hbo9mcYHFNQLAdGMHgBYMSvqAQZ0U1/wsPBCaEFsO30JDa/DjfMjJVUX0ZjF
Mez8w0t2s7xP67juPkv2lmHSb59HeXu8sMtGqX1LYpyXnAmwTTGHoHolE8pHP1tGv3ebAstOlQMT
3bASLp0MIWtwdjGPWdryM91QVCcDHerp+Zqc8rIbnbNW7wz7kr27dRZ/3NVkGdObk5M+LfJEk2KH
9+F+UZAeZiyLlesMDfeVuj4rcyY8H+xMH1fZN3h196u7lYa+WoJV0L1wv+6b92nIEnWf/wQsQ4Oa
k+B4QuLlEq3FWmEqwRdLjC5HYWmzs2sP9O/okQXh7AiZP+U4FDCpNTDqJYwCAmPoPJ5F16RSNbhj
gRAXA9bHAOeClCiqdbU0cQEzPI1AopNA+NroUHFRiGeV439720erN9OX6ZwCPxboPkz9o6UaJ1qH
f3ndZgJh26oFxeQKk8nF+LCKM4iYwsUvwKYoIkXT3IdJDSlUviT+NIPZRU9nOqdiVSlj0hy6RYEC
ad4fsIAd1Bah2JdnhSNLS3/SzfKl6kf09C724iZJ+Lve5uDBZwUGpXsspd8L2YmOnsXj0okTHQq+
t37mlHsohgXqwnrlKdm+H2w0v55D0oHj7M8L0UqHPHm8WrO0l0vF6MF41u2CLxms/es0apadziWE
zjwlX9jjI7NzOpKiJT8cZTq9h1Iaw8UYyU3bn+43UmZvns7jNRWUL9K5RYiPf4x7FAy+UhChiS5O
EjeDDUn10Ntq1h5gZen3adKgDU2KFsfk9WndPbCEUR/uNBsOZsbjs11X1nr1YobJNKuo1eMs1PbH
KN1EC6kJL9ii0oXESTnovPh57S24hDy0oAV//DJK7SRZDbZh8zsynQPxSstNlh2eYPJ/JOx2e18k
WTzVF13wfu1PmxKLo3Y5vLP1MjRPHG5S1TCndv16WVtAC9xZPsFdwE97pdX7t8vis7Zq9ABWDM3Z
C+um8jHiE28HiuPAbaAmA25VdT4/SYushrDryd2LaYM7fbgIF7JHJBR0IqfdjBYeC4HbI5ieTTvY
1iPyfX6CE8YCIG2LcG8jOi7zCySZbiNPY2pxXyhs4SEMrX24LKNCv5mxtZl5neyBk3Jc1bOhP4lr
ZlNYa7lkbdGoeQusz3R1QExU65figGrRbwMzbAQQ4dQeA/DQAYwsbby47T1kOH4m58aGhx1FbHQq
qAikFENlyfa47mMRbhWAGKZMZlmdWTsN7UIMEB/qnbmbWGvl49PD6o+DzTRiJk8kQuxFH5Pygclh
gvbrD3xojhMc0zZJ4Iseqhv1ScG4GAquXXpWXB078xmzdPsVWHqZG78p8GM94OcBJHOy3R/PDQl7
H1UIFZfu9do4jNN/vP73JKmmygi1/y8IALXstf7OeKxbZkPV9H3aLnh3kRKsruOvIoq10M1ew8ZS
KWLOg82vM6PpJ1BCLVdIU28XZ4A4xNBYJv0EsVP5WQxAR86Sw5vCk3ppvDSFavmHWAL3ZvC7lrkv
MuhmvXs/xy371vNVvClByJiBdxxC8MsYGDV4uu5yxuPG4k4EaXPwZsPjM9fWcyXUWY0lBp7rBJjE
HTnmIUBbwD0FVrxTKJXvlpB/B1xRNSW8DGq5AimvDzuGh0yKeo7kTjk9JIXj4KbQiHLZjRv+yl4t
3itYjz/9tx0LjyRUZiAFO7loMJz+RAY4KGG9slep60GI2S+OCFosOnnZbFVqhTWJy5b2FO14BoxI
+jTXhuPhNQ7Y//sYrRQhHV3MilKR4MwQlrk8OLAEwU5GgXHeCX+8ItMoaWCJu3AFtvmqBhfRV0o9
j840PDEra7R8acY0KIvHi9Lu2jlWwJPEU+rgvjj1luT+rqYUu+pTsi3rBCenWjOLLakotyoV+sW9
Dtml5sDaOfMio+EN50eTRPGysLmF/ajpDtfeGbg/KEwsLNjsMOdJHIouiKdg7Zpvvsqy9mqHu+c/
2WO8Asht8gqEDkbeCnqiqTX5HU8HbYnS1Ba3JoMANp97PZ+wMp9sopYf99Yw3KmW0owhOOBIOsnF
RcYLiZqgZS2/HEzIrvoVpuNu21AtOe2/3R6FbKwRzK7pFl8ZOL3fzMcCBJZG7KwDkirrp7Vi7Ars
i4tQAp7Y/RkSVJslybMlwLnXAFzVh/TDizSU8K3WeYBQx44PvPGEPuf9alt6ausBg3Ib4vUmNG+4
HDCtUHKBx0ncQDn5cJUx8kej28LGHjDJirUpv3bdnFO+m2ogtygCI2rYJC0mNxxqNvIgQRWdLwfK
lXnVUUE2gKj7zZ3g4P9OBQvLtfCDbssveQw4M4283X6ryN6ajqIu5/EKxnEjKjgB2tG4TqCPrIsR
qZOE97j9VLtCxmqrhbEAxO1hdXppy9x4WO4sgHKQRf0E1RTIf3K2eT8c85hmm71pCGLPHDtbDC22
vz8yRGrYq9U6n2eEIEt3resepuoubrq9+FCcHdFBYrHSwlC9aZtnRdt10TTx1mvX187SEUAQ5RnL
wDFJgZE2zVbuhCGxhusd5PTTW3GBPERANF1+P3vJHUEFJ44lJNwzXKtuf227aBRPq7IwpMsdi7Vb
TwhFBOccrgpLMR9eR/SOBPOJTrGXEjShwQGgS/Xcnc/lTN4asjL5kORF0cwmwoJ8lXmjPCgoydrn
L9v8lLuzJJ/LJNxiGqD6q/Kaxq0yRrKgFFSk/ul+WfRrCgBhlil5/6OvSm3BqOy1JxUVV2CeylHA
dcYXQcQC3U582cb7d1j4tY4iXjFRL+hzvicPZODTGQCtnl/br09Kj6F8fMWaWaTOiPcdtUfsfUjM
X19dL8EeaxOBA9Nqsi0Kbel4Ehm2qJJmG/Lw15zy+SOri/EShOwEusx6VEyh9I3e6w93bo405QU8
5SI6EgfWU8DdXrQMdv78SlIR141ihVDSiuDjhTehp+24ML95Hh3/4GaCFy/mLJEInw5kkQ/BtKh3
aHaVYIOs66piLS6aU40qJ7l7cYjWeo/ZAerZMFe775/auPxoH6fOmuZcjboVKWeW99agckMEIpjS
RS26cQUZkKg2LQEuZCVk4U6TNnmr4W0cz+rZdetuSoiWFxCpeWlh4v7qwrim5tHAnqEr9HqJab0P
MBI75I72KVDwOGqHYqz5/fUCMVhyi8ngEy5bAi2A1MX9h5AE5UlUfteUBV44hA00jBsq6qM4ZWEc
ez1HpNj6rZwfsBUtuSaNRa6rcEk/6olOD4Pj7mLU84q3S5g1SUoX6JmyHa0pl7EpKeKZzd+gI6gI
cxLitClKbcvsyv9zUA/U86ZgNl/YsCO2Jq7O9iSHQkIrW6Rm7/RZb/bIuB9QWSIH8ynjbC2GZDHN
PSTUoFqbWxaq4jnaFjmZV4wc5F79n0PhGTeF22P0AjVQzHXtQW6GyG9/kN0Asd3MDcWuYi9tQQT7
OzKuXcoLbZaJKZxRzAtr0ViWBLKvYWTUCfrPIrJuETE6/dK2G9XRup5mL+Qp5ZTYrQK1RvpvVBLu
fZR3yZkfN7k+pWMQrAUjJDBeg7bUsZyjV85qkS8GDR1sbwgWlAQIJaZ3dmSY0BIAFj9y/4H75yzN
Y9egBHQjXwmw8zp0GtsctvrEvHbSDMjyBoM5GmAIUZ3oaUNy0HMXphfBxLngMMuqOH9oAc2ypsdi
QNApYif44aDibyCZ8qrflYqka3cXtL3SAFCWXXWWPgxd+Rq+DlluzK1opSkAqmiUtIGG73BzpHOu
515w1Gt8gj+6H5HnCEDOlNH67Ri61pXBQLu1iDwpYUpV9VifZCZ+V1EM32YNuMqRSvDbeVfxhCvP
jRrWt9nVcSL7Lp2AMPpnNDi9/4zxLufKrxSg2+uLxltP9aooddxGgTrNEyHDI3OBD2PhsKDKKVom
0rd4M3cXYucOwtuYm8UXISc+UZ0jFtOz9mAtE5Oex45Bil+Lk2Wuw4UG1MypbW3S5eJFgl1Qhf/+
Jxl6aQp99vN01YyOCP53mPN5WUxNVeLMpha6BgD6Y3GDf2ynPQ6AcerLv48w8UP8j/G1H5VwkYxb
Coxhx05aok4vqetYUI0kvJTMaM/qAbMQUmRYkRyCU85Rsg6DifZcz+U4t4m6XpUUJRLhwZ7vpTeL
p6x7+mNzNCVOQvNa45bx4nRm+QuAtuaK0k9enMllVlzqrMz0HucUVOvJ1lZgeDLyFH4cXO0bcY/Q
iqEcN0RxUFZ1Rb7xhC6xSxOBpZ3k7MzOxLbqFodtOYV0RYGeOkFE4Fqx1vxOeyx5eVYLLLRPf5K7
Rxa62Fj/+r7L47Dc7XFLB8wgYTeKzFLZPetwU3XlZRAJ8MCBU5/bojWS5oVVQ2X9YkcDqsCEHVy+
++SESGjaYv8M5gy5tHpFshaNgSVo5sTXuT9r177uCZUFub6Kk1is55caH2J4RZ0Owbn4qkNC+g23
L4e7GEyqa6gX+oVxT7dx/KyJW8TU7NDdHf7fwuae75h9Y/VyWl/O7C14+3JJmsCiDv+ovGzuONw6
SfJqSNf6ohFwkbOSMXHZG57w63bJZbU3H7SDvp7UWY7hd7FrVWmJZpEJdmat3s//VwUGegXHcKjl
ZJjXO2RhhPcvIF+JyCv9q0CnlYTCWuqMtdHmjkC5ga6e8Q6AMQ28bc+OssV6HR6Dx/x4NUH2/yKy
+zrdGJIudwuT532pBrpVzLOSWH7PCbrdK7tLn0jq6NYfmRbersN7ic4GlDe/UiEY+DrS5VtCTUa1
hFTb7qGgV3NbFAOza8witoPUjXtdTJ8HpPKXPATpPLfA+hyRZ1TL5dSPFIjOWBdZcu5zLr7f46nX
5WYHduu8FD0hJY5QxcB9cOUVfazXQwF2Swlhm/AwmDjD/2IHcX6nDb612TNZHW46XQCzb6zcFcTe
uk4xPqF+UXu80H5fo6BhyJl8pxzLi55+GQ7EI5ZeXSX+uAJbtmhgvaq1Q3+PuARezzY0aomIaYjS
iSgbfnRWLuV5spU/oUaeXeSSIcaFeWPpe10dPY2jN0o2ACosR99ztRzsDjNoafyrK9fwUbzA6Kfl
9dFsYl44mlB3EGHvSn3Y8RiojZGxRy+xvQfKitoHHIDdBWL9xLZvclLSjWgXehFYPCNJ3mn1Wgw4
StjtXWT7c+d2vKQHM5UiYD8Fljo97o/WRxQ0U/xirH2R5CEaCeO2bjg6MEc5HpNKMWXbE2L9ccon
Xu+4XFhKssrq/pU2navSKS2b9JsyeS7phjTEfFV02ZWO13uUUTgvMoISTBysyVGJsU6S/eetMmOm
HupjxlWbEqcRdEJTlusTbX2APAJ163nh1RaKv/WJnvhJ/jglcBRG+1FzaYXQhajkSf3uzHorO6dI
HkBRVAgfBLdCT8ovOIESCZYhezljeLqVO37FiL+OZR4TAS/tiSc1g4DSdUD0Epg1ZYA7lZYfBPQ7
1iYFsl3iRv1gRwqnHOfKAgmxlWa0MOZeC8pA/GtKbCH2hRRzBB7nAWWRVMZQRGspRd1N2JJgNJCX
AwPJ1Jw02ggMOWVmeGkKM32gx8qp1YTqV4HIe0szuuYjMHbGTATXYIZ1r0qI8GCoyDU1bKdAiYB9
HQGPO47jkUQGAyFQbZ/9eJ8zJMQrc56mPi1HZz1+v7YzBl2wD3Moghg/1xIxSxtGK0QZHh+VZN3z
Ji39moFTNOpaT9+KcJCw8KhNGGiUkOPOXJACIrp8w+/O9Hzm96y1v7bv+VhbUo5fRnN6f2jKTXY9
IaAkFSZxOw3wCTP6S/vtwjtet/z9++geuopw2avO/z/OIVuex2NWXZ+Nbh5bkU/hnbE48D18QCh3
Do/y9OTIrIcUWG5EwI0pJLbbDnso3YtEIi/Qy4DJlbI8tTeZOnm92l2pVevtwe1BXjRwx2aDo/Sz
kclvWXZoI4ymzW6f0GWxKHvWjxvpLAZZeLYmIWmU5/33nt08SEOxAKbUP+x41dSk3LesUSpu8+GG
I4RXflXI9nxgmnAMkvn//WfLVvM1zPKdXf9qpWune39xl62K44kqJZrBKGBIAzYafKhQ6/QzYltK
rLWy6XUpPiEWYIbKTYz1yIib1IU3rCbnPmieDBo92s44YRvaP/cVVSjIyQ7rQQSEfcC+UVHkjUSK
uzGU9nBrHAcsb7tgXiZ6OI/QTpWLPbp6OEUl9JljXwSMhXzwGA5gcHC9h6J+bp8pOoZa+QAZZRvz
ZxGT4QuHFSDz/KnXJDBtaQvEIahQ1ecy3LnIKn/w0DjWPYdNP6TJnC/v4ONvmHuS06V9wuArDoZk
f97/2O4i6VMGzLhBlRBo/w11ZcXa6vfQk4930c2N/Eo93IksueYCmVSAAKtvxwDlQr1GIXGTHKij
tHtde+TW+PG9x9PWcPdAtgr86KUVBeGo+ztwz/NhtCAkYePbe+5YpuMxzhOPwZreC2162d6J+PHa
uzsypGkuRAcYFprlYgEYXHNND7qi4It3XjauLWxcpOCyXKJBAv72VuIr/qQ1fEiGAdyVMpDWM/la
J9aG4i5okTwQfE7ksQ1MDD6DDRkNCsts7JF8+PNkLPX9va9kunMXPOuH2v1xvBIyM75Clizxcdzs
aZxBZncGYWycPGNVjEhSZ95u8UxGfqHWCgvaKPmPObzYgeBY5Q42+vjpcGNkMM5aqT4bOiowoAOj
nAHUHSGg6ZpoDVI2c47nR6j8cq7ToUjd/GaiMRiVjXKAHNwuuKSYRbqGwK42wEroy0zJblIgsaCu
m3FwG2myw0oHp95i9t1wnsPl3VREQLA5/iHEwAbLbxNX5WVh5TFXsflyG4VY7ONAxozRPiAaxTEl
mhj4R4Hq6vzhmcfuG9DXNuaP86BlyUVNJsJguhP17N4bMvspCFZ5nOT+avBxe6S4R9HUbmvi94Ss
rwlCIwVVf53KOIvnz7Rfj687+yE5t/ik+2Geo/UbEJhT/M3iBPP3LG6IUamL3dR0FrJrDnpSUu1I
XVxA+XRx7l/G/mcIP9fwyFzJGW80vIyNlNsYy5HzD8cJEa03CuzUH/ivf8U8QCPFrC6GzSvdZlSB
f+y4aRb0Bs/xY/SIxbA4yaFxaV7VHsI+k/kBHiJsBGqOSkbK6ixH4J08489DiZIp2NOFCxg/IQzt
QOknIBbvZzTFdSA36E8lkxgLhItOxSwm1gslJRgarTsOwbl/+ySKf31PsS8idMCF3+OR5Ne1L9Ax
UlRBU7MhHzlgSHuoUmAc8z52sF0Pd5SYeCpgpkJy1v3i6EaEW3VQhVgNyBacaDwfr/Oo3KEZsWnF
Gr70K8oafiDqDVxL1BlAVYVRqyv+3t++4THP1UDyuGz7Les9Jn/ZiT3ewneO7IxD1yZ5Rih1CJ4c
6l0lDtbglAP5BGlZr4BnLWIdnBiXKpaTlim4QvJWRW5xDKtz0KV5DI+ICtLp9MrX0271pnUZ6xky
raTLAz6Laqbo7OpC6bZ18ucdvLAU4LmnDRKyF/TXd6UMcaeEY3C3o0zLBx+UWrbltHSTuN8Ie/jJ
n5Qp4cyVMOTEP4JXNmUDabLJroZCgmceVVNJuP/rpeDJcblLMMTbXCpMDWvUBBlYXhmk4Nq1sCEd
W5YQOI95wtJ3lTPm4UqaAek4E6eo5RmQt7Y0l9zkxuNoT0jhP2SiLIFqS83bzESNnzapG4WWbRcQ
hEiVpFe/ze8dTTi4ruRnO+/Cxjk5CweIDPKm0toxxIuIhVhPww0pxsoODb9ZVuUMInh/zZmJ+03U
tDQcIRyZRE2xEkmXOOdp380DHz1DSPw3g8saTmy7UJ940QwyjTg8MCoBzE8iRYpGdxE0CLYAf0w9
fkvYRPxHh1Y6ndJEM+nXh7gLW7qvEqXBCumQ10MfCqlRYGYMZmuF3gxpO1BOs/UWQtNn7fPRaZcs
nX5I3udvV0lwxG7pM3txva8f/KiL/Sii4plzy8KdXMuNyZETEhH4td+exmCtLFePo7B//MRG/g8H
4ToA5ud1gAKRPKIPDkW5/a5hboZYPLz2x+vlM5vSkMBnrcPLXl8T8UuI7f43mV2NYwwGV+gLejBQ
0KmeMmQaRktgjYWbu2eGw1Qm9hFdwqzFo37R7dO9flbezj6nm2l3QPAOYUsJ2iBCWpyrFJMvAR30
cywSvvlAaoIMwIVpTzUmaHgpYET5hOGK5nHuQha+4XPokxTL6Y00dyOb4Ls7srmhC8SkhRMjOeo7
9h+iu1EUGumlehDvjEb1k/9ndwqViDtX34k8uF+inLLQ4n9g+eX3KMQ59i5yKhyB50mZ+TBOi5CC
AKCuNd18KFpaYLdTmviT6d40rlbb2KCus6xbh5h2tWX8d+1KWhKM1H+VWy0uRgpM5etk9Z4MLBi4
dSLwmVCSS0PAaWbCLikm97C97X/vG5mMl9vsqzxkB0PXBH8TgJBAlfcBlL6xqiCGp71zNUYW+sXr
fp4TURcqIocYZDBdLRVd/7InQ4u8/CqYmtqwgH1kDGhh3MhXKu148Zyqm7Djsyhs5x/HJZWmAm/1
/Z1h4rhwjmx1GQf4OSL/v0t1kx15XMBbj3P6oz4ndhahyE4lA5u5s6uQyltlgGUVrU3WWoDuaBHN
Gf0iqHWVspm4N2owD+4mGuqxoqSl80kbF86H/n2xHvk4i8XKoUsccLmfymMLQxnMb649Eefp6HwJ
1fE2WPiWBvTOr5D9rXKzz4fS687P4L40or03fU2iqqJXGovGX8ZAyRnO80Sxy65CBpHjUMUvIqNw
fZHGEZOw+ijNSRDjLqF4lE5lj4dJNiZLFuVRbYOvZPWTJL8t7lAJBrb/DGGEzgyr+i3mFuyJk2JV
sy8GIAkBT5k2FchxX36VohWaKFS5MFzqfxYj2iI9sfDquk6+UtCGzBqncWHCWq75EPJH6lhpewNy
F9Ed9xJsMlGS0ZmlfCI51bgSyDSBXQUdu1m2F2qk9rACRdua3U6p0CzFcvIqeB3vwy4srjRma3xg
lbtgSPxjJYm99axkSgrojZo+t/R024UQ/YkVml6xuKNP+qhEceZZ87KNA14uY/eRsl5mTHmjzMCl
oVrlcU09Pr0ynpty/2vXh6LeGz21fmLOHa3XUDhGGWRCUmfvCrLG06JwDk8s4CaCEj85tQuRAtGZ
UiiQqdgQr9wRvIoV/QWgKNVyQiBUIm48aNlp7hSMestuoBnX6Vqv+aUnyCRuRh0JdiQcqnkuNCoL
XRT18PHLNBgpAdbjEXMovBy4kkJTy/sCblmnV+vPbeJh0hG/XxqSwiDJESuTv7Et7Dyo0zSaT7qI
1QPUVl/yRZijVwYI+d9jLOPcnOkgYMLPiOqcHIEMyC1wEZQHJIaFyuoyY22qF124pM3OsApbahd1
/Js1H+AcX4jUSYUEcIfTM/P/54XUpSvgsw5xoXbi9FzoREy0ExWD66/RS69V1mU8JfMoCgInowf7
dJsy/f2b+DyQSrGQxji0RaN+jNHGyxGdLbrJLcFRLM1w7EMM96vKLBmO0zpk5LnLWFzyk0sqsKgS
Vn+Fe6sRzHaDVis/bVZLnQ0uW71KvUaTdThi9LUxpuD0MpSg+DbDWlVfvFYsU6ulyBSBgvM0Qpgq
/YjzcIStRoGvM8YP2kf/58jRiDnJCV7xIqXEes4FCppEtrw5jx79sySk2MccFOX+p3ekhraSAdDj
9Riax0H3UA7veQyi7rLknm+Wq7DH5Au1BjGdvXTVQ/KuIf5luQBdMqF7Qu8XN8DFFzkru2KJR2DY
2Ex3bdlYgiy0JImGBN2d+ZGmHD4sJLn06XW/9hWQmE0zDvdc+DJbpw27GjOLYc0PH1c2/uRtTrad
oL44SnCOeiuIu3u3EkxN73lUWC1pWBQrcHFtddH6NEVQcq5xA+LwCbv2o0j9CDvNAv6Ib0z5wbTt
l1nAJFtWvupf63ZlDM9xTo6cOGLD5zvJ0HNpVlOWHwTs7CETO9tAnL4fZrgVo4B7Tw+6+2HzRzzl
Q8VyQA7xIXs3qDT2k+2gqem5kJy72C209qzieZiwVWyGtSnCBF022m7+hJuPaVFeVHtei9BrKV5W
fGlTOlHWGX4RN0+2dKgdFG7cShPLJ3BVnxX8Gjm4kY8mKmhJ2dUKPyZfLNxyzGTigK/45gumY5k/
6+FHm6QdkBQOe1HvRAr5ZwCjdt+qy7QXxPXhrwLZD89r7KE+doJS76/QIy1h6HGxVc0nd2I+mGUI
Qr46ZeTNugzWnkDKCD+AGyDh+GqazaVgGQ7rMqsDE8S4ZQREfPUe/PnyjoUkDc7HZwhF0YruEVsR
A56vqRiLhcXs1/n3wXjpVS9ANru59k50WHypaIDod2Ebe1wWXFvqCtMnX9tbyXi/fRm2fm99YQJo
nElF1c3OMvy0esl9+efCcLDRYBYCwTj8iSxJX2Ic4RaltMK8F8YrLQVUfZMuXugyLzee36+Akzs9
MyyryKtC1BT74C7I2xho4i57YxXze+H8KRjp+V2LoWXlVPqmzZNTnu/9RSeZGawSBYq0MpoEZEaN
TQ1bgTcPFMMtD6N+xL+9rb71+IRZgA3T5eAxFE4ol3bnZLSORK4pbC1tZIKDtRDlVh1aWimCX8/S
1LgOGsVfJNWIUPssUz9rH+1QHuIAh3hrjz7z75jzk3K1b2DVCWANG2yF0v6k72v5j339R3zkdJzM
eMBiCK/8G6oBOMtGCnmF1EkvXlx1LKogt3ZrZkQLv8S+zHYCxsOg/CyhgfExFHtbz7zun9XCJn36
xnYhDJTZNcyS355lUDY063SpFZmr2hOXRF2rwTfuOCrbOhmy6Mn8cjnPKUc2zgaeq4uxw8Uti6ih
wd46sIgKJsYXvD6LzIpB9mPaHjRw3bMzmUkWtDOzAfTq9Yx8I6p/CE1L5gHNtiqbi1jfatz6PioE
y6YszmPniCdit+1xKQRLjUKAXVFtaYqRF4yVY8iKorUFZSY9goGDdbGltu3FSmG7CIqD+m0dga4y
BBocb+8ZX1XPt/R1MXin/DaSngdglGALI7KoFgT2VJwdLJUx4MRbRiams7oHok4aQSl33FAXfzJt
ELvf1Dj6HIuTvxUYmokhGYrO4SBHk5REFYrs+zNayI5FMCreAMHUNGOG9etDMJULjsKg2bZwhXwp
Ww16oEeTbboptC+njdBouK60vvLcU98DyXY+6VszmU3psGH//q2Cw1/fN9UeKnAd7cfcx181jyBm
WtH1c0WdEGa+gh0zaBIO7SUXuqHONgTGsEbbguAftGNC+HMBbtI2Au5NFruV70vqjK3wihNOaToQ
VqtDz8ZA4XTa4JNNsmHaynf8WGPSt0G9WANTynuk3S3KkASGE5B8QOAJO6Ju4UiXj7Co3U5SSnlU
ygkkdtZyeo9FeVrjdOtS4m4jG/FK4Js7PY+MFVqLMdZV2G6QCyYMSsb4igPo6lO8Xx8i0cs6SSio
4Xl8GTrsfdcD2rCJgp+irqa6kzTBewwunvJvy0hFYWq04lngRfxA3uc7cY96DmJma/5/2xFmf/fS
56+n4ovnWLCrf4kzV5DlwDRK/zhhA/rFAPwyrZ0YV6ZTkXlgHGX+Pz6iuV59tRSpLo+hGCofYQ30
yImJXsGkBYa55iBjQZ90ekjStq7uaxjHl8zIh4nYU1HrX2Mw5NR1LzMfqsYaf4bHAeqWKqnehxIb
TYwfaXs0hVyU90kuDKU1D2I1rzbZtl4Zy/hnJ36RSrtPhfVFL7BaPfwX+9A2g1z1sJ9ooR/rj1y3
In0CmTf+/WMJ1GSZj7kO0wrLsHK+qFAxtfCpRI5HCuJvktMXru6soKbs5+iXJ9k8ODof97kjkmMK
oo+eVCObAFJCx1FRaSCbj1zF7rYsE6j3CmCFapQ5crzGTAF+dAgiIgt/ADZFP/ygveLFAC/O/n3r
9m6I+7/6Xg5dUaUlCnysr7BxQ1Uc4D+MfgzkeWt17lwj94DZJTS3QPuw/36mB2xKg+KHsrVcdE7I
s6G7E1pB73/vAoca/3cacB4RKMEvZalJ/SmrIqV1WZkqV4KwutP2DZC1SHKe/cU0RUZH/oBaig7K
7IvxKcp/lYb71p9QD8JxvA0p8Jj1Ps6GG+zA61r0lhKocJnyp9Ync+Hnjs9jvQ5XYiYI8FhmWHxq
5MiHFACwMZAJKM2/UzSw/+IuuJ3FesaCK9ctl7O9iVvMKlPuCv7z8hQ95m9kpInGk7hLO2i1sRFk
YTAJOUiRhmEbiAPm2hNatgM26/ekEQuS9eJxDeWegsYsqnUQZVHu1ts/XX3QnaMWaqregZhLANoi
5IsRPJQ0ZX7Gyjp2PRdjnftTWxwl/Y+zKj1YKCKIdX6vQhBKl7snxgLdSMMBr5A3RpJFYasnDsIo
3VNv0oU/riUocPZBq/VEg/DNjfHCH5ePxYNZVNOgC0XpF183mBx5gZO/LLNp9BNC9Gbc9GUz/9Z0
2SL6oXVAAfJJpvO8dtIJyUxfUY6cuvbLKC5XX1hAcg4L7i/0p1w2ipRj3rFiUNJp0oqKnpXYhJ7u
YG0gInZCQJRqfFYqpAXLkV8WXxyJUjtRS+svzjFqggFtbjo3iB680ufkeC8OXtvDKatRxw/Y5qSk
se8p1CZ/hZ+qH6RyNw2QZ/X/Z/u/nndmPJNCTWgRDbxjs+nQKDQvtdoixU3ORR3qkbSoRd9QYp/l
PnpYh7bOLGsuX5tLyp5YN8okzZJOAQVyF+RgYZo3NyLpIzm9aSz9LNRWqTrwmyFRf1JlenXvFFYf
/UVJDLKHlet7Yqp0Fho9Og9DL61s8lYOMHTmEq8+LkgsI1Bmom0fe0CASMejTnN0WRJDJMcJHgEz
qtSHRTGZhTjmO8TxcZWrUQShl/rfcbD+hrqYhOHpBv/8GPi8AFqh+rIhmPfHU8j11k0dN0Ljzqjq
O5GxPaCXebOiQgvVcL3WAff3jqJQeNY20JDdIbGkxBosFABH2zG+h2s830oxA4UV9J3KIZSjvDZl
oHHzEKzwh4w8iDMCTl4DUJMQT44JhyLrktbP4QWR323RIqqzP/UAXW2qqXD8o0ft0UP+fCo0rQoG
92IHKjwhacV+zCO3K0D/RV8gxSpQWXId8PlIIu1Jws9DsHa1lLQCylQyzM+wY97UCW1O6m0A0nqc
c9tco5eGvfcBhy+flbB0k7cZlH1SeWk34O6MsoIyinP/qldFOjDhQjIV4GFMyp8JUpd2o2bkO3x/
PrmVGImITD7YO1Os87cg56XvceoRzndTmvsb2zH1TFLf6x4h/pd4LkHh2lHPoT3an6ziQXvPHxe3
nPLk89HqWRwE4x/eeS9S7jFWiF7sx8f3lFjHG6qHnQhnQF8lY8Af9sIBEGv3EyDZpCsY7/KrjuOt
lRHtbL99FTWT9xEG5tQZ0AAUug2jThMJW37j1m1fdo8gugDGBaze7T6ZOxHRnk9kixBfokvC1dOS
JBoFkowoIRMBfVdjY5kuaHo3JAwMlAFnHxKGK+fkyy2dVN1dlkjqQiO/qJ2IoBODZapY6+CXn19m
U6/XHgIgO5KE7e9lSKtGf5nxAnv96bZAOXir8iuS6+l/Xppp+C8Aqeid0Wq0HYC1zWpVhigMa3CM
oXHVwt0VHIn4sXKTr+EWuZGdyO+CTcBNJRwndSzahZn2nGKgy3MzSd9El4fjJyWmxF1KGxNwDqpQ
AoWG3bkRTTpRlybC6qyvBGxhOvoGHZUE9cWqTlzuTSFuXE5dixj04XXoNWSBy8SLITFauSzMotgx
0A6JpjKlUB9NjlQXIwdbymz0aVgs0BFqWdLB9IfhdzpVSiKmRIATsb6gVDtKREEjZdBaaD78nQU+
vpt90sLLLev7PKQ8utbtnaxF5Qs6GA9xaYeBOXE/EzNptPWuxZ/9OT9s7BGop1zQK8Xn5mYy6v0Q
7Efg9UNszmK+ty+ofncKMwiWJkr2eZkzKscg121dMtulbTOXORnBOZcjKtNf72V00pKO6Sl0k8xy
qgW+iIPegz6kPIKQkD5J0g8TYJY9VwLSK2aFQE279g9q4r1lv4maV5WBgewoTBxsTd0dURZMtUz/
kSLBViffONFyLkwhIgkxkYeNIkPU7xJuZsDbQ9ttYieeRfqQmc5bWEe6Ja1q2bOTHMb23lB8OKuU
vZG5OfxmwTMVMbAz9IaPu9v8p7nvYPUTk3YIixpd6d0X6l+BqBlTT9PQM1r+Zu2YPHABDnejgFyN
IezWjo/YcAwGlxdKOy5mryyTL7uOOR/xC5YEP6XL6MfcFaE8nGTWwtZAw+NDkSLceDjxHdDksdoZ
PLZr72jMmxWREbm1uUIaVjAVNgxWYeaYlAq5LRFoPDaPHr6s3kUo2CrA1esJ39r12BUes6Nn9Nza
rVT/wUJj5V6Tq40AiZWBB8wqcc3EMkgV/HOXgGkXdiGK78mQ7004qcA45rVxn02JigoyWiWZmweK
BsFEfYjZvIf5TBpRpWlK/dpxcQZ2vpNPYR3MXdHZQkK57mK5bKhYjcqTNqWudqMS8VFOFpZUjvFE
u9EunOy+cFsf7Gf9QoFQmLGpsxsANRDT+SjBe8Wp/q1CBBX39k/wITWaWTyANGHvCloEMQSspmqQ
tQWQyirhuuSrumdcU9oM3o41io/StrWGN/7uoe6X5RShHowtsLF6RNnfUICciCYwFfBtyN+siqm6
U9N+0w8EkdKk5uUbO5hcrCldfPFFDx1cTJ0T+wIO3Wwfvi7vOBfmqBs1+d/JAD+VN5EyCjJtWnZK
NYDk05+5/im/5I6BRWwje3TW+kQYwVsEIqjCemfCDhWnkf/5rKuw5XVoOzB0IVG8u3RD1enfD5vX
HDoxxgm9T8CWWo755ydA/CfB68qYqNA7VycnSZBA545E78QBCRJC/tP9ni5faNMZMnRkf0TI82vn
mjnWx3wgFzC1xPWqra7fMPeiEzf/JSaBi8zIa4padbHdMgGAEJI5OxsQ5wcgN4wE9Vzu9mjtp+Dj
ZhBwvf0vgIRyKIcfm4KZsp7be+/t8UHMIkcOl84RBTbo2b3WROyZthHUQ1g37M4lOAUMaw0WzFFh
ZirFU7cac5cSdXlrDSK0KLZSz7ldNFINvb53ZdrXXAvbb5WotLrMcE2ct4x3lWt3zvs3z6MStjC0
5KiKToyLpB8W1r8Mg/ZBV1FB14e5mcsPR6w0yeuefJTEJ2xQo9mSbNZLgelQ6nTzcpQ/hBWHREBq
2Ovd729YWYLzRN39xzBXDAu/l4GHqiCyMxJAYUW+zZkgyxUEdoEAPQAv4SNHjBPQY7hSBPRDyFO4
msSL1oVaD+63GVhFFFCUC7XKNfIfQQL9k+N3HIg3rvD+lkdnMTIxPSX1HSdPQUCglDlvFjtjys35
M0HEaSxjAZz2s3yRQaJR7BGkk3VRiq21CMgKJqfKlClWr/23Z0lpfK1epLVbeTqaD9nDNLqAAdkf
SByZBjp1f1zrRiksHZFNxUxbH7NjKHVwqrlWtLLHlEfw7Bt5BmMge2skDaPsR5ISn2Fz+1YKVDSX
BjUlyVlkpANw9y3peb0IMiG6qjkpLrMSAJp+OJE871ExUSkpoZQLj80NHklnLuHxD3Emf/1BM9Hr
FaWb1jooHMMlcULZf7nJagG+jhncp2myARJ3aElV0eRv0aD/RqiOEec69m/kGEB5Zw8VA1RKif4O
beyPCa5wNhF0kt5AwJdg5BKksfc1vMksVOo6c1gUafoLSJ1jLTEtceU/Nc/WECKtpRcg/hJF/qXu
cAQ67hPHQg0iOd5hGWRTKdYcBZegY4asO8Ng5Ukq8ojfhcV6mpQmDmoBQ6UXUYltEdjwUCnNlgMt
pid5TaObn9h8GWBEQMmiMQPnNl3/WhEEU5AwfcPhTRHF98DOOaN5fn8eTeFSWtVSnAzC2pV1cB1u
tGcs/9m69UIJCE88Unrhw2fk99BvggqTErIelUcvzTtiMqvV3TjfehZaAtHji4rtqodcFlovnRK7
GuO9GunAws2cxQH1vQTHIozziCUvabdMydNVwf7SADk7dyS6BaJ9jH1Tq+tgkxvBXXVUFtr0evvk
CpeOUiy8BohWB727oD8je27QUotjubMXwFL/qNoymQJvyD+uwLo3nE1I0xA0AJvaZuqh4OKlo4te
i6O7rt9f2VIxaTE3AyPATtJoMFYjZiKXyiqVWqhpkOVz9yfH9zvNGI++rE/uEOeP51PYtMqkRnPL
cEdEwO0Qh5kz7MYv5IHLvu4lJn9B5ChMVK9XJ0GfLZoCQvMBpqNXFNG1V2ePa98suLhYVAi2WnhW
q93OpuvlUgilbawPmX/DgXlJF1RZkC9VBvQYBC+nkgJTOiD70/4l/gbj1p1glHPiEKVaQ68pS2kZ
JnKoUsoTCA5CqYOsFR/+76OLA/IsW3Fw4cp+uvN5D9hBCBXBjGxIlKWCOaV3OWfXokLp4cLHdAX/
xdIOfgfVz5taKcsz+dW3AKJXTlugecwhgCOwlZM2DQJ50Pf7Dnee3OoHMp2PxmAdBojpFVgjpwkz
y7vHaTB6q6O9FhoIyhKhBRiFOy+UwzZSTHYntvcOqLFfWrgGUFMETxiD/bxAXX1cgcxqesaQOpLj
ytccnml5221SZK555Y9dR9AGDlbB/340e+n4S94YlmPW6rohVhw9E+WjlVfah6OVHYfThv1eBP7A
CzaJkSTqUUQAN7hkMP2qKoNo3agEPGVwcOKv7hJrCVNwQmZZCc+sQiNd1LfP6/ysCFHcPd9BwIii
ZtGxxd5NQ8RV9DuLycNZgnpPhbI56MnlQBc9kqXxzbgWiX6MXhm96pJxiyF3RkNaYQYaPn+nGV4v
7Uc3O8MgVuiAvZxMeycLuQNKFUEyi1x4Dw9QGScSR/pN8VdoEJNhs7qsft5V4WCZzwoICLOXWOhP
vj6GiR4iebJcI7mIapMuhht5wVRH9o2woCQo2ao32AHvBFehweGuO6vaUbeFnBqSgP1j0MyVBK2X
gcwsq+doFhHqgQWJSTTmj5w3vCf3yC69bfHZygdqhyR+71JL+34KwZZ2sZRKu1rshKE2hSly291H
LEh7y2mRubVJc1zNz5JhxbfbgiJdUs1Eqgw3sqfyFfozpr/tc8G2J3jWuu3CGIFcf6rtFiAT0n8q
VuPwzi226/7vXm8ge9padfhlCAGdbh0AuCydsflYnq0lrQVrAmeq0ebTfrNrSitcZJ3i1rMcvntN
POquV9QOtVeoJxb1+C3cr04pZnttuK+fa8HyxOaj2KfIlWM3j78ooSgihpa8y6oXkFgkXhQkeAmN
yYIpzw4lKRSU6q9KV8oA8ESxu8ABya+XNn7teRZ6WciudK7eCsKZLeTa3QJk79En5pmw6Rt1mYP1
jJhgPf4dut0buvV5g2F8TsmzIJm7KWG22qcKdgVAAH14y7sTSlbpDpy0/QzXmw+l9aCHRMNkIbdo
Q5sOAC6X/OvYmM5xKku9PtYRsbMHoxtU3OKLHC0ecXY0Ll8sVFcW84OjHtjWy7WHyq0PYL61wUQ8
yPg/vp9v5EbpSmhmyct9S8gij9reFcwKOSihT7K6B+VtSSUHeco7lnCGsGg6ytkn/c5uwOgRzVco
yjbdKRTFn5/FBXM1gP/zm30T/sh/p/ZEue4/6ymtMqIPEB+wfaG2K1+60NyevztdoQM8vDgFbyNF
Ro9oQ2ck/8UoY6aV3oxGspsnyn9093Kn1F5QGkVsACq2Fhv8UGm6vTeko66T3geKtsRG4ds+RarM
DftyKIpj7IIIj7+moU9QPuf4GsKltuHfVmzHMrsekbd2q1QNARMvs+gmCtXI5K1qUZb5aEGi00U6
eiga9WeAN9uYXxnIi71DY2oZ8NAB0vm0CqUIz1C93jhKsLYnTc8Fr6E5PomTRGlYCjWYCV1WmbjK
CM67e3yOo22mbmmzzQTuy07+rxwsINc8dUCHa79cX4lz8bT++0EsNlZnHtW+OHIjqKWHsR3+QOQ1
V5VFYxMr/JLVW1keMXunYs/vjf2ODerYga2zW3vF5dAzeuWF4JnEz+SoNIfO8/I4wWhmiH0BbV+h
eWJoI0vd3de4vNtDuAamW9ol3D6Ot+FdlkbptgM/mXXNFAH3IGLESAqrooTXN0nMXzpcklxHgmO0
2+myXO7Os5lntpbwMW5J1LHZ0DWS4/oSk91b9zkL0TgQutb2WNDYzaQ31BTfMeqFU9x5qLoX89CT
sWhbKbthf4bRrh5sYL0XsNwGb0/4bmbotS01YuTnLiusVKAt5aeOWXYL9zH1pB94
`pragma protect end_protected
